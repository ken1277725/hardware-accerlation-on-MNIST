


module recog(
	input clk,
	input rst,
	input wire [7:0] rx_in,
	input wire rx_valid,
	output wire [3:0] out_number,
	output wire [2:0] out_state,
	output reg number_valid
);
	parameter int = 25;
    
    wire rval;
	onepulse ONP (rx_valid,rval,clk);
	reg signed [int-1:0] NN [0:7839];

	// DFFs
	reg [783:0] alldata,next_alldata;
	reg [9:0] alldatapos,next_alldatapos;
	reg [3:0] number,next_number;
	reg [4:0] pos,next_pos;
	reg [2:0] state,next_state;
	reg [3:0] anspos,next_anspos;
	reg signed [int-1:0] max,next_max;
	reg signed [int-1:0] ans [0:9];
	reg signed [int-1:0] next_ans [0:9];
	reg next_number_valid;

	assign out_number = number;
	assign out_state = state;

	parameter GET_DATA = 1;
	parameter MUL = 3;
	parameter FIND_MAX = 5;
	parameter FIN = 7;

	wire [391:0] data_in;
	assign data_in = (pos[0] == 0) ? alldata[391:0]:alldata[783:392];

	always @(posedge clk or posedge rst) begin
		if (rst) begin
			alldata <= 0;
			alldatapos <= 0;
			number <= 0;
			pos <= 0;
			state <= GET_DATA;
			anspos <= 0;
			max <= 0;
			ans[0] <= 0;ans[1] <= 0;ans[2] <= 0;ans[3] <= 0;ans[4] <= 0;
			ans[5] <= 0;ans[6] <= 0;ans[7] <= 0;ans[8] <= 0;ans[9] <= 0;
			number_valid <=0;
		end else begin
			alldata <= next_alldata;
			alldatapos <= next_alldatapos;
			number <= next_number;
			pos <= next_pos;
			state <= next_state;
			anspos <= next_anspos;
			max <= next_max;
			ans[0] <= next_ans[0];ans[1] <= next_ans[1];ans[2] <= next_ans[2];ans[3] <= next_ans[3];ans[4] <= next_ans[4];
			ans[5] <= next_ans[5];ans[6] <= next_ans[6];ans[7] <= next_ans[7];ans[8] <= next_ans[8];ans[9] <= next_ans[9];
			number_valid <= next_number_valid;
		    
		end
	end

	always @(*) begin
		next_alldata = alldata;
		next_alldatapos = alldatapos;
		next_number = number;
		next_pos = pos;
		next_state = state;
		next_anspos = anspos;
		next_max = max;
		next_ans[0] = ans[0];next_ans[1] = ans[1];next_ans[2] = ans[2];next_ans[3] = ans[3];next_ans[4] = ans[4];
		next_ans[5] = ans[5];next_ans[6] = ans[6];next_ans[7] = ans[7];next_ans[8] = ans[8];next_ans[9] = ans[9];
		next_number_valid = number_valid;


		case(state)
			GET_DATA:begin
				if(rval && alldatapos < 784)begin
					{next_alldata[alldatapos],
					next_alldata[alldatapos+1],
					next_alldata[alldatapos+2],
					next_alldata[alldatapos+3],
					next_alldata[alldatapos+4],
					next_alldata[alldatapos+5],
					next_alldata[alldatapos+6],
					next_alldata[alldatapos+7]} = rx_in;
					
					next_number_valid = 0;
					next_alldatapos = alldatapos + 8;
				end
				if(alldatapos >= 784)begin
					next_state = MUL;
				end
			end

			MUL:begin
				next_pos = pos + 1;
				next_ans[anspos] = ans[anspos] + adder;

				if(pos[0] == 1)begin
					next_anspos = anspos + 1;
				end
				if(pos == 19)begin
					next_number = 0;
					next_pos = 0;
					next_state = FIND_MAX;
					next_anspos = 0;
					next_max = 25'b1000000000000000000000000;
				end
			end

			FIND_MAX:begin
				if(ans[anspos] > max)begin
					next_max = ans[anspos];
					next_number = anspos;
				end
				next_anspos = anspos + 1;
				if(anspos == 9)begin
					next_number_valid = 1;
					next_state = FIN;
				end
			end

			FIN:begin
				next_alldata = 0;
				next_alldatapos = 0;
				next_pos = 0;
				next_state = GET_DATA;
				next_anspos = 0;
				next_max = 0;
				next_ans[0] = 0;next_ans[1] = 0;next_ans[2] = 0;next_ans[3] = 0;next_ans[4] = 0;
				next_ans[5] = 0;next_ans[6] = 0;next_ans[7] = 0;next_ans[8] = 0;next_ans[9] = 0;
				next_number_valid = 1;
			end

		endcase
	end


	wire [int-1:0] adder;
	assign adder = 
				(data_in[  0] ? NN[  0] : 0 ) +
				(data_in[  1] ? NN[  1] : 0 ) +
				(data_in[  2] ? NN[  2] : 0 ) +
				(data_in[  3] ? NN[  3] : 0 ) +
				(data_in[  4] ? NN[  4] : 0 ) +
				(data_in[  5] ? NN[  5] : 0 ) +
				(data_in[  6] ? NN[  6] : 0 ) +
				(data_in[  7] ? NN[  7] : 0 ) +
				(data_in[  8] ? NN[  8] : 0 ) +
				(data_in[  9] ? NN[  9] : 0 ) +
				(data_in[ 10] ? NN[ 10] : 0 ) +
				(data_in[ 11] ? NN[ 11] : 0 ) +
				(data_in[ 12] ? NN[ 12] : 0 ) +
				(data_in[ 13] ? NN[ 13] : 0 ) +
				(data_in[ 14] ? NN[ 14] : 0 ) +
				(data_in[ 15] ? NN[ 15] : 0 ) +
				(data_in[ 16] ? NN[ 16] : 0 ) +
				(data_in[ 17] ? NN[ 17] : 0 ) +
				(data_in[ 18] ? NN[ 18] : 0 ) +
				(data_in[ 19] ? NN[ 19] : 0 ) +
				(data_in[ 20] ? NN[ 20] : 0 ) +
				(data_in[ 21] ? NN[ 21] : 0 ) +
				(data_in[ 22] ? NN[ 22] : 0 ) +
				(data_in[ 23] ? NN[ 23] : 0 ) +
				(data_in[ 24] ? NN[ 24] : 0 ) +
				(data_in[ 25] ? NN[ 25] : 0 ) +
				(data_in[ 26] ? NN[ 26] : 0 ) +
				(data_in[ 27] ? NN[ 27] : 0 ) +
				(data_in[ 28] ? NN[ 28] : 0 ) +
				(data_in[ 29] ? NN[ 29] : 0 ) +
				(data_in[ 30] ? NN[ 30] : 0 ) +
				(data_in[ 31] ? NN[ 31] : 0 ) +
				(data_in[ 32] ? NN[ 32] : 0 ) +
				(data_in[ 33] ? NN[ 33] : 0 ) +
				(data_in[ 34] ? NN[ 34] : 0 ) +
				(data_in[ 35] ? NN[ 35] : 0 ) +
				(data_in[ 36] ? NN[ 36] : 0 ) +
				(data_in[ 37] ? NN[ 37] : 0 ) +
				(data_in[ 38] ? NN[ 38] : 0 ) +
				(data_in[ 39] ? NN[ 39] : 0 ) +
				(data_in[ 40] ? NN[ 40] : 0 ) +
				(data_in[ 41] ? NN[ 41] : 0 ) +
				(data_in[ 42] ? NN[ 42] : 0 ) +
				(data_in[ 43] ? NN[ 43] : 0 ) +
				(data_in[ 44] ? NN[ 44] : 0 ) +
				(data_in[ 45] ? NN[ 45] : 0 ) +
				(data_in[ 46] ? NN[ 46] : 0 ) +
				(data_in[ 47] ? NN[ 47] : 0 ) +
				(data_in[ 48] ? NN[ 48] : 0 ) +
				(data_in[ 49] ? NN[ 49] : 0 ) +
				(data_in[ 50] ? NN[ 50] : 0 ) +
				(data_in[ 51] ? NN[ 51] : 0 ) +
				(data_in[ 52] ? NN[ 52] : 0 ) +
				(data_in[ 53] ? NN[ 53] : 0 ) +
				(data_in[ 54] ? NN[ 54] : 0 ) +
				(data_in[ 55] ? NN[ 55] : 0 ) +
				(data_in[ 56] ? NN[ 56] : 0 ) +
				(data_in[ 57] ? NN[ 57] : 0 ) +
				(data_in[ 58] ? NN[ 58] : 0 ) +
				(data_in[ 59] ? NN[ 59] : 0 ) +
				(data_in[ 60] ? NN[ 60] : 0 ) +
				(data_in[ 61] ? NN[ 61] : 0 ) +
				(data_in[ 62] ? NN[ 62] : 0 ) +
				(data_in[ 63] ? NN[ 63] : 0 ) +
				(data_in[ 64] ? NN[ 64] : 0 ) +
				(data_in[ 65] ? NN[ 65] : 0 ) +
				(data_in[ 66] ? NN[ 66] : 0 ) +
				(data_in[ 67] ? NN[ 67] : 0 ) +
				(data_in[ 68] ? NN[ 68] : 0 ) +
				(data_in[ 69] ? NN[ 69] : 0 ) +
				(data_in[ 70] ? NN[ 70] : 0 ) +
				(data_in[ 71] ? NN[ 71] : 0 ) +
				(data_in[ 72] ? NN[ 72] : 0 ) +
				(data_in[ 73] ? NN[ 73] : 0 ) +
				(data_in[ 74] ? NN[ 74] : 0 ) +
				(data_in[ 75] ? NN[ 75] : 0 ) +
				(data_in[ 76] ? NN[ 76] : 0 ) +
				(data_in[ 77] ? NN[ 77] : 0 ) +
				(data_in[ 78] ? NN[ 78] : 0 ) +
				(data_in[ 79] ? NN[ 79] : 0 ) +
				(data_in[ 80] ? NN[ 80] : 0 ) +
				(data_in[ 81] ? NN[ 81] : 0 ) +
				(data_in[ 82] ? NN[ 82] : 0 ) +
				(data_in[ 83] ? NN[ 83] : 0 ) +
				(data_in[ 84] ? NN[ 84] : 0 ) +
				(data_in[ 85] ? NN[ 85] : 0 ) +
				(data_in[ 86] ? NN[ 86] : 0 ) +
				(data_in[ 87] ? NN[ 87] : 0 ) +
				(data_in[ 88] ? NN[ 88] : 0 ) +
				(data_in[ 89] ? NN[ 89] : 0 ) +
				(data_in[ 90] ? NN[ 90] : 0 ) +
				(data_in[ 91] ? NN[ 91] : 0 ) +
				(data_in[ 92] ? NN[ 92] : 0 ) +
				(data_in[ 93] ? NN[ 93] : 0 ) +
				(data_in[ 94] ? NN[ 94] : 0 ) +
				(data_in[ 95] ? NN[ 95] : 0 ) +
				(data_in[ 96] ? NN[ 96] : 0 ) +
				(data_in[ 97] ? NN[ 97] : 0 ) +
				(data_in[ 98] ? NN[ 98] : 0 ) +
				(data_in[ 99] ? NN[ 99] : 0 ) +
				(data_in[100] ? NN[100] : 0 ) +
				(data_in[101] ? NN[101] : 0 ) +
				(data_in[102] ? NN[102] : 0 ) +
				(data_in[103] ? NN[103] : 0 ) +
				(data_in[104] ? NN[104] : 0 ) +
				(data_in[105] ? NN[105] : 0 ) +
				(data_in[106] ? NN[106] : 0 ) +
				(data_in[107] ? NN[107] : 0 ) +
				(data_in[108] ? NN[108] : 0 ) +
				(data_in[109] ? NN[109] : 0 ) +
				(data_in[110] ? NN[110] : 0 ) +
				(data_in[111] ? NN[111] : 0 ) +
				(data_in[112] ? NN[112] : 0 ) +
				(data_in[113] ? NN[113] : 0 ) +
				(data_in[114] ? NN[114] : 0 ) +
				(data_in[115] ? NN[115] : 0 ) +
				(data_in[116] ? NN[116] : 0 ) +
				(data_in[117] ? NN[117] : 0 ) +
				(data_in[118] ? NN[118] : 0 ) +
				(data_in[119] ? NN[119] : 0 ) +
				(data_in[120] ? NN[120] : 0 ) +
				(data_in[121] ? NN[121] : 0 ) +
				(data_in[122] ? NN[122] : 0 ) +
				(data_in[123] ? NN[123] : 0 ) +
				(data_in[124] ? NN[124] : 0 ) +
				(data_in[125] ? NN[125] : 0 ) +
				(data_in[126] ? NN[126] : 0 ) +
				(data_in[127] ? NN[127] : 0 ) +
				(data_in[128] ? NN[128] : 0 ) +
				(data_in[129] ? NN[129] : 0 ) +
				(data_in[130] ? NN[130] : 0 ) +
				(data_in[131] ? NN[131] : 0 ) +
				(data_in[132] ? NN[132] : 0 ) +
				(data_in[133] ? NN[133] : 0 ) +
				(data_in[134] ? NN[134] : 0 ) +
				(data_in[135] ? NN[135] : 0 ) +
				(data_in[136] ? NN[136] : 0 ) +
				(data_in[137] ? NN[137] : 0 ) +
				(data_in[138] ? NN[138] : 0 ) +
				(data_in[139] ? NN[139] : 0 ) +
				(data_in[140] ? NN[140] : 0 ) +
				(data_in[141] ? NN[141] : 0 ) +
				(data_in[142] ? NN[142] : 0 ) +
				(data_in[143] ? NN[143] : 0 ) +
				(data_in[144] ? NN[144] : 0 ) +
				(data_in[145] ? NN[145] : 0 ) +
				(data_in[146] ? NN[146] : 0 ) +
				(data_in[147] ? NN[147] : 0 ) +
				(data_in[148] ? NN[148] : 0 ) +
				(data_in[149] ? NN[149] : 0 ) +
				(data_in[150] ? NN[150] : 0 ) +
				(data_in[151] ? NN[151] : 0 ) +
				(data_in[152] ? NN[152] : 0 ) +
				(data_in[153] ? NN[153] : 0 ) +
				(data_in[154] ? NN[154] : 0 ) +
				(data_in[155] ? NN[155] : 0 ) +
				(data_in[156] ? NN[156] : 0 ) +
				(data_in[157] ? NN[157] : 0 ) +
				(data_in[158] ? NN[158] : 0 ) +
				(data_in[159] ? NN[159] : 0 ) +
				(data_in[160] ? NN[160] : 0 ) +
				(data_in[161] ? NN[161] : 0 ) +
				(data_in[162] ? NN[162] : 0 ) +
				(data_in[163] ? NN[163] : 0 ) +
				(data_in[164] ? NN[164] : 0 ) +
				(data_in[165] ? NN[165] : 0 ) +
				(data_in[166] ? NN[166] : 0 ) +
				(data_in[167] ? NN[167] : 0 ) +
				(data_in[168] ? NN[168] : 0 ) +
				(data_in[169] ? NN[169] : 0 ) +
				(data_in[170] ? NN[170] : 0 ) +
				(data_in[171] ? NN[171] : 0 ) +
				(data_in[172] ? NN[172] : 0 ) +
				(data_in[173] ? NN[173] : 0 ) +
				(data_in[174] ? NN[174] : 0 ) +
				(data_in[175] ? NN[175] : 0 ) +
				(data_in[176] ? NN[176] : 0 ) +
				(data_in[177] ? NN[177] : 0 ) +
				(data_in[178] ? NN[178] : 0 ) +
				(data_in[179] ? NN[179] : 0 ) +
				(data_in[180] ? NN[180] : 0 ) +
				(data_in[181] ? NN[181] : 0 ) +
				(data_in[182] ? NN[182] : 0 ) +
				(data_in[183] ? NN[183] : 0 ) +
				(data_in[184] ? NN[184] : 0 ) +
				(data_in[185] ? NN[185] : 0 ) +
				(data_in[186] ? NN[186] : 0 ) +
				(data_in[187] ? NN[187] : 0 ) +
				(data_in[188] ? NN[188] : 0 ) +
				(data_in[189] ? NN[189] : 0 ) +
				(data_in[190] ? NN[190] : 0 ) +
				(data_in[191] ? NN[191] : 0 ) +
				(data_in[192] ? NN[192] : 0 ) +
				(data_in[193] ? NN[193] : 0 ) +
				(data_in[194] ? NN[194] : 0 ) +
				(data_in[195] ? NN[195] : 0 ) +
				(data_in[196] ? NN[196] : 0 ) +
				(data_in[197] ? NN[197] : 0 ) +
				(data_in[198] ? NN[198] : 0 ) +
				(data_in[199] ? NN[199] : 0 ) +
				(data_in[200] ? NN[200] : 0 ) +
				(data_in[201] ? NN[201] : 0 ) +
				(data_in[202] ? NN[202] : 0 ) +
				(data_in[203] ? NN[203] : 0 ) +
				(data_in[204] ? NN[204] : 0 ) +
				(data_in[205] ? NN[205] : 0 ) +
				(data_in[206] ? NN[206] : 0 ) +
				(data_in[207] ? NN[207] : 0 ) +
				(data_in[208] ? NN[208] : 0 ) +
				(data_in[209] ? NN[209] : 0 ) +
				(data_in[210] ? NN[210] : 0 ) +
				(data_in[211] ? NN[211] : 0 ) +
				(data_in[212] ? NN[212] : 0 ) +
				(data_in[213] ? NN[213] : 0 ) +
				(data_in[214] ? NN[214] : 0 ) +
				(data_in[215] ? NN[215] : 0 ) +
				(data_in[216] ? NN[216] : 0 ) +
				(data_in[217] ? NN[217] : 0 ) +
				(data_in[218] ? NN[218] : 0 ) +
				(data_in[219] ? NN[219] : 0 ) +
				(data_in[220] ? NN[220] : 0 ) +
				(data_in[221] ? NN[221] : 0 ) +
				(data_in[222] ? NN[222] : 0 ) +
				(data_in[223] ? NN[223] : 0 ) +
				(data_in[224] ? NN[224] : 0 ) +
				(data_in[225] ? NN[225] : 0 ) +
				(data_in[226] ? NN[226] : 0 ) +
				(data_in[227] ? NN[227] : 0 ) +
				(data_in[228] ? NN[228] : 0 ) +
				(data_in[229] ? NN[229] : 0 ) +
				(data_in[230] ? NN[230] : 0 ) +
				(data_in[231] ? NN[231] : 0 ) +
				(data_in[232] ? NN[232] : 0 ) +
				(data_in[233] ? NN[233] : 0 ) +
				(data_in[234] ? NN[234] : 0 ) +
				(data_in[235] ? NN[235] : 0 ) +
				(data_in[236] ? NN[236] : 0 ) +
				(data_in[237] ? NN[237] : 0 ) +
				(data_in[238] ? NN[238] : 0 ) +
				(data_in[239] ? NN[239] : 0 ) +
				(data_in[240] ? NN[240] : 0 ) +
				(data_in[241] ? NN[241] : 0 ) +
				(data_in[242] ? NN[242] : 0 ) +
				(data_in[243] ? NN[243] : 0 ) +
				(data_in[244] ? NN[244] : 0 ) +
				(data_in[245] ? NN[245] : 0 ) +
				(data_in[246] ? NN[246] : 0 ) +
				(data_in[247] ? NN[247] : 0 ) +
				(data_in[248] ? NN[248] : 0 ) +
				(data_in[249] ? NN[249] : 0 ) +
				(data_in[250] ? NN[250] : 0 ) +
				(data_in[251] ? NN[251] : 0 ) +
				(data_in[252] ? NN[252] : 0 ) +
				(data_in[253] ? NN[253] : 0 ) +
				(data_in[254] ? NN[254] : 0 ) +
				(data_in[255] ? NN[255] : 0 ) +
				(data_in[256] ? NN[256] : 0 ) +
				(data_in[257] ? NN[257] : 0 ) +
				(data_in[258] ? NN[258] : 0 ) +
				(data_in[259] ? NN[259] : 0 ) +
				(data_in[260] ? NN[260] : 0 ) +
				(data_in[261] ? NN[261] : 0 ) +
				(data_in[262] ? NN[262] : 0 ) +
				(data_in[263] ? NN[263] : 0 ) +
				(data_in[264] ? NN[264] : 0 ) +
				(data_in[265] ? NN[265] : 0 ) +
				(data_in[266] ? NN[266] : 0 ) +
				(data_in[267] ? NN[267] : 0 ) +
				(data_in[268] ? NN[268] : 0 ) +
				(data_in[269] ? NN[269] : 0 ) +
				(data_in[270] ? NN[270] : 0 ) +
				(data_in[271] ? NN[271] : 0 ) +
				(data_in[272] ? NN[272] : 0 ) +
				(data_in[273] ? NN[273] : 0 ) +
				(data_in[274] ? NN[274] : 0 ) +
				(data_in[275] ? NN[275] : 0 ) +
				(data_in[276] ? NN[276] : 0 ) +
				(data_in[277] ? NN[277] : 0 ) +
				(data_in[278] ? NN[278] : 0 ) +
				(data_in[279] ? NN[279] : 0 ) +
				(data_in[280] ? NN[280] : 0 ) +
				(data_in[281] ? NN[281] : 0 ) +
				(data_in[282] ? NN[282] : 0 ) +
				(data_in[283] ? NN[283] : 0 ) +
				(data_in[284] ? NN[284] : 0 ) +
				(data_in[285] ? NN[285] : 0 ) +
				(data_in[286] ? NN[286] : 0 ) +
				(data_in[287] ? NN[287] : 0 ) +
				(data_in[288] ? NN[288] : 0 ) +
				(data_in[289] ? NN[289] : 0 ) +
				(data_in[290] ? NN[290] : 0 ) +
				(data_in[291] ? NN[291] : 0 ) +
				(data_in[292] ? NN[292] : 0 ) +
				(data_in[293] ? NN[293] : 0 ) +
				(data_in[294] ? NN[294] : 0 ) +
				(data_in[295] ? NN[295] : 0 ) +
				(data_in[296] ? NN[296] : 0 ) +
				(data_in[297] ? NN[297] : 0 ) +
				(data_in[298] ? NN[298] : 0 ) +
				(data_in[299] ? NN[299] : 0 ) +
				(data_in[300] ? NN[300] : 0 ) +
				(data_in[301] ? NN[301] : 0 ) +
				(data_in[302] ? NN[302] : 0 ) +
				(data_in[303] ? NN[303] : 0 ) +
				(data_in[304] ? NN[304] : 0 ) +
				(data_in[305] ? NN[305] : 0 ) +
				(data_in[306] ? NN[306] : 0 ) +
				(data_in[307] ? NN[307] : 0 ) +
				(data_in[308] ? NN[308] : 0 ) +
				(data_in[309] ? NN[309] : 0 ) +
				(data_in[310] ? NN[310] : 0 ) +
				(data_in[311] ? NN[311] : 0 ) +
				(data_in[312] ? NN[312] : 0 ) +
				(data_in[313] ? NN[313] : 0 ) +
				(data_in[314] ? NN[314] : 0 ) +
				(data_in[315] ? NN[315] : 0 ) +
				(data_in[316] ? NN[316] : 0 ) +
				(data_in[317] ? NN[317] : 0 ) +
				(data_in[318] ? NN[318] : 0 ) +
				(data_in[319] ? NN[319] : 0 ) +
				(data_in[320] ? NN[320] : 0 ) +
				(data_in[321] ? NN[321] : 0 ) +
				(data_in[322] ? NN[322] : 0 ) +
				(data_in[323] ? NN[323] : 0 ) +
				(data_in[324] ? NN[324] : 0 ) +
				(data_in[325] ? NN[325] : 0 ) +
				(data_in[326] ? NN[326] : 0 ) +
				(data_in[327] ? NN[327] : 0 ) +
				(data_in[328] ? NN[328] : 0 ) +
				(data_in[329] ? NN[329] : 0 ) +
				(data_in[330] ? NN[330] : 0 ) +
				(data_in[331] ? NN[331] : 0 ) +
				(data_in[332] ? NN[332] : 0 ) +
				(data_in[333] ? NN[333] : 0 ) +
				(data_in[334] ? NN[334] : 0 ) +
				(data_in[335] ? NN[335] : 0 ) +
				(data_in[336] ? NN[336] : 0 ) +
				(data_in[337] ? NN[337] : 0 ) +
				(data_in[338] ? NN[338] : 0 ) +
				(data_in[339] ? NN[339] : 0 ) +
				(data_in[340] ? NN[340] : 0 ) +
				(data_in[341] ? NN[341] : 0 ) +
				(data_in[342] ? NN[342] : 0 ) +
				(data_in[343] ? NN[343] : 0 ) +
				(data_in[344] ? NN[344] : 0 ) +
				(data_in[345] ? NN[345] : 0 ) +
				(data_in[346] ? NN[346] : 0 ) +
				(data_in[347] ? NN[347] : 0 ) +
				(data_in[348] ? NN[348] : 0 ) +
				(data_in[349] ? NN[349] : 0 ) +
				(data_in[350] ? NN[350] : 0 ) +
				(data_in[351] ? NN[351] : 0 ) +
				(data_in[352] ? NN[352] : 0 ) +
				(data_in[353] ? NN[353] : 0 ) +
				(data_in[354] ? NN[354] : 0 ) +
				(data_in[355] ? NN[355] : 0 ) +
				(data_in[356] ? NN[356] : 0 ) +
				(data_in[357] ? NN[357] : 0 ) +
				(data_in[358] ? NN[358] : 0 ) +
				(data_in[359] ? NN[359] : 0 ) +
				(data_in[360] ? NN[360] : 0 ) +
				(data_in[361] ? NN[361] : 0 ) +
				(data_in[362] ? NN[362] : 0 ) +
				(data_in[363] ? NN[363] : 0 ) +
				(data_in[364] ? NN[364] : 0 ) +
				(data_in[365] ? NN[365] : 0 ) +
				(data_in[366] ? NN[366] : 0 ) +
				(data_in[367] ? NN[367] : 0 ) +
				(data_in[368] ? NN[368] : 0 ) +
				(data_in[369] ? NN[369] : 0 ) +
				(data_in[370] ? NN[370] : 0 ) +
				(data_in[371] ? NN[371] : 0 ) +
				(data_in[372] ? NN[372] : 0 ) +
				(data_in[373] ? NN[373] : 0 ) +
				(data_in[374] ? NN[374] : 0 ) +
				(data_in[375] ? NN[375] : 0 ) +
				(data_in[376] ? NN[376] : 0 ) +
				(data_in[377] ? NN[377] : 0 ) +
				(data_in[378] ? NN[378] : 0 ) +
				(data_in[379] ? NN[379] : 0 ) +
				(data_in[380] ? NN[380] : 0 ) +
				(data_in[381] ? NN[381] : 0 ) +
				(data_in[382] ? NN[382] : 0 ) +
				(data_in[383] ? NN[383] : 0 ) +
				(data_in[384] ? NN[384] : 0 ) +
				(data_in[385] ? NN[385] : 0 ) +
				(data_in[386] ? NN[386] : 0 ) +
				(data_in[387] ? NN[387] : 0 ) +
				(data_in[388] ? NN[388] : 0 ) +
				(data_in[389] ? NN[389] : 0 ) +
				(data_in[390] ? NN[390] : 0 ) +
				(data_in[391] ? NN[391] : 0 );



	always @(*) begin
		case(pos)
			0:begin
            NN[0]=25'd0;
            NN[1]=25'd0;
            NN[2]=25'd0;
            NN[3]=25'd0;
            NN[4]=25'd0;
            NN[5]=25'd0;
            NN[6]=25'd0;
            NN[7]=25'd0;
            NN[8]=25'd0;
            NN[9]=25'd0;
            NN[10]=25'd0;
            NN[11]=25'd0;
            NN[12]=25'd0;
            NN[13]=25'd0;
            NN[14]=25'd0;
            NN[15]=25'd0;
            NN[16]=25'd0;
            NN[17]=25'd0;
            NN[18]=25'd0;
            NN[19]=25'd0;
            NN[20]=25'd0;
            NN[21]=25'd0;
            NN[22]=25'd0;
            NN[23]=25'd0;
            NN[24]=25'd0;
            NN[25]=25'd0;
            NN[26]=25'd0;
            NN[27]=25'd0;
            NN[28]=25'd0;
            NN[29]=25'd0;
            NN[30]=25'd0;
            NN[31]=25'd0;
            NN[32]=25'd0;
            NN[33]=25'd0;
            NN[34]=25'd0;
            NN[35]=-25'd1;
            NN[36]=-25'd5;
            NN[37]=-25'd29;
            NN[38]=-25'd178;
            NN[39]=25'd304;
            NN[40]=25'd697;
            NN[41]=25'd268;
            NN[42]=-25'd61;
            NN[43]=25'd260;
            NN[44]=25'd780;
            NN[45]=25'd346;
            NN[46]=-25'd44;
            NN[47]=-25'd40;
            NN[48]=-25'd28;
            NN[49]=-25'd10;
            NN[50]=-25'd2;
            NN[51]=25'd0;
            NN[52]=25'd0;
            NN[53]=25'd0;
            NN[54]=25'd0;
            NN[55]=25'd0;
            NN[56]=25'd0;
            NN[57]=25'd0;
            NN[58]=25'd0;
            NN[59]=25'd35;
            NN[60]=25'd13;
            NN[61]=-25'd10;
            NN[62]=-25'd164;
            NN[63]=-25'd207;
            NN[64]=-25'd416;
            NN[65]=-25'd839;
            NN[66]=-25'd994;
            NN[67]=-25'd1162;
            NN[68]=-25'd1485;
            NN[69]=-25'd1853;
            NN[70]=-25'd3109;
            NN[71]=-25'd3843;
            NN[72]=-25'd3421;
            NN[73]=-25'd2918;
            NN[74]=-25'd2099;
            NN[75]=-25'd1629;
            NN[76]=-25'd1075;
            NN[77]=-25'd699;
            NN[78]=-25'd420;
            NN[79]=-25'd132;
            NN[80]=-25'd13;
            NN[81]=25'd0;
            NN[82]=25'd0;
            NN[83]=25'd0;
            NN[84]=25'd0;
            NN[85]=25'd0;
            NN[86]=25'd0;
            NN[87]=25'd78;
            NN[88]=-25'd78;
            NN[89]=-25'd963;
            NN[90]=-25'd1330;
            NN[91]=-25'd1659;
            NN[92]=-25'd708;
            NN[93]=-25'd1667;
            NN[94]=-25'd2274;
            NN[95]=-25'd2075;
            NN[96]=-25'd3790;
            NN[97]=-25'd3235;
            NN[98]=-25'd4758;
            NN[99]=-25'd6434;
            NN[100]=-25'd6692;
            NN[101]=-25'd7127;
            NN[102]=-25'd9137;
            NN[103]=-25'd9594;
            NN[104]=-25'd7307;
            NN[105]=-25'd5458;
            NN[106]=-25'd3766;
            NN[107]=-25'd1750;
            NN[108]=-25'd685;
            NN[109]=-25'd156;
            NN[110]=-25'd35;
            NN[111]=25'd0;
            NN[112]=25'd0;
            NN[113]=25'd0;
            NN[114]=-25'd3;
            NN[115]=-25'd9;
            NN[116]=-25'd134;
            NN[117]=-25'd1670;
            NN[118]=-25'd2373;
            NN[119]=-25'd2088;
            NN[120]=-25'd1697;
            NN[121]=-25'd985;
            NN[122]=-25'd2521;
            NN[123]=-25'd1780;
            NN[124]=-25'd5202;
            NN[125]=-25'd3035;
            NN[126]=-25'd4299;
            NN[127]=-25'd2341;
            NN[128]=-25'd4947;
            NN[129]=-25'd4129;
            NN[130]=-25'd6256;
            NN[131]=-25'd7218;
            NN[132]=-25'd6154;
            NN[133]=-25'd6697;
            NN[134]=-25'd4714;
            NN[135]=-25'd4551;
            NN[136]=-25'd4182;
            NN[137]=-25'd1326;
            NN[138]=-25'd214;
            NN[139]=-25'd4;
            NN[140]=25'd0;
            NN[141]=25'd0;
            NN[142]=-25'd13;
            NN[143]=-25'd93;
            NN[144]=-25'd655;
            NN[145]=-25'd3158;
            NN[146]=-25'd3741;
            NN[147]=-25'd4643;
            NN[148]=-25'd4212;
            NN[149]=-25'd3735;
            NN[150]=25'd268;
            NN[151]=25'd871;
            NN[152]=25'd1095;
            NN[153]=25'd9139;
            NN[154]=25'd11955;
            NN[155]=25'd13925;
            NN[156]=25'd14416;
            NN[157]=25'd18832;
            NN[158]=25'd15365;
            NN[159]=25'd5363;
            NN[160]=-25'd204;
            NN[161]=-25'd232;
            NN[162]=-25'd1860;
            NN[163]=-25'd7414;
            NN[164]=-25'd7734;
            NN[165]=-25'd3428;
            NN[166]=-25'd923;
            NN[167]=-25'd197;
            NN[168]=25'd0;
            NN[169]=25'd0;
            NN[170]=-25'd10;
            NN[171]=-25'd177;
            NN[172]=-25'd1253;
            NN[173]=-25'd3185;
            NN[174]=-25'd4712;
            NN[175]=-25'd5697;
            NN[176]=-25'd6451;
            NN[177]=-25'd8825;
            NN[178]=-25'd2842;
            NN[179]=25'd1082;
            NN[180]=25'd2955;
            NN[181]=25'd10887;
            NN[182]=25'd12978;
            NN[183]=25'd11289;
            NN[184]=25'd15035;
            NN[185]=25'd20472;
            NN[186]=25'd21410;
            NN[187]=25'd12788;
            NN[188]=25'd9510;
            NN[189]=25'd11258;
            NN[190]=25'd9122;
            NN[191]=-25'd3141;
            NN[192]=-25'd12797;
            NN[193]=-25'd8134;
            NN[194]=-25'd3070;
            NN[195]=-25'd503;
            NN[196]=25'd0;
            NN[197]=-25'd9;
            NN[198]=-25'd123;
            NN[199]=-25'd599;
            NN[200]=-25'd2566;
            NN[201]=-25'd3657;
            NN[202]=-25'd4776;
            NN[203]=-25'd6845;
            NN[204]=-25'd10694;
            NN[205]=-25'd4622;
            NN[206]=25'd266;
            NN[207]=25'd5714;
            NN[208]=25'd5714;
            NN[209]=25'd8548;
            NN[210]=25'd8905;
            NN[211]=25'd9840;
            NN[212]=25'd13613;
            NN[213]=25'd21248;
            NN[214]=25'd21150;
            NN[215]=25'd14796;
            NN[216]=25'd8233;
            NN[217]=25'd9553;
            NN[218]=25'd11632;
            NN[219]=25'd5421;
            NN[220]=-25'd8644;
            NN[221]=-25'd9566;
            NN[222]=-25'd3527;
            NN[223]=-25'd18;
            NN[224]=25'd102;
            NN[225]=-25'd46;
            NN[226]=-25'd317;
            NN[227]=-25'd862;
            NN[228]=-25'd4097;
            NN[229]=-25'd5868;
            NN[230]=-25'd6049;
            NN[231]=-25'd7767;
            NN[232]=-25'd7210;
            NN[233]=25'd439;
            NN[234]=25'd1802;
            NN[235]=25'd3430;
            NN[236]=25'd7697;
            NN[237]=25'd5349;
            NN[238]=25'd9724;
            NN[239]=25'd15795;
            NN[240]=25'd25431;
            NN[241]=25'd22786;
            NN[242]=25'd18038;
            NN[243]=25'd11801;
            NN[244]=25'd8753;
            NN[245]=25'd6197;
            NN[246]=25'd15039;
            NN[247]=25'd16254;
            NN[248]=-25'd2548;
            NN[249]=-25'd9637;
            NN[250]=-25'd2873;
            NN[251]=-25'd120;
            NN[252]=25'd0;
            NN[253]=-25'd14;
            NN[254]=-25'd218;
            NN[255]=-25'd769;
            NN[256]=-25'd3931;
            NN[257]=-25'd5788;
            NN[258]=-25'd7403;
            NN[259]=-25'd8018;
            NN[260]=-25'd6511;
            NN[261]=-25'd553;
            NN[262]=25'd3951;
            NN[263]=-25'd168;
            NN[264]=25'd4462;
            NN[265]=25'd11299;
            NN[266]=25'd7741;
            NN[267]=25'd4847;
            NN[268]=25'd16055;
            NN[269]=25'd22640;
            NN[270]=25'd21727;
            NN[271]=25'd17277;
            NN[272]=25'd8760;
            NN[273]=25'd3008;
            NN[274]=25'd12690;
            NN[275]=25'd23041;
            NN[276]=25'd5059;
            NN[277]=-25'd9046;
            NN[278]=-25'd2893;
            NN[279]=-25'd67;
            NN[280]=25'd0;
            NN[281]=-25'd15;
            NN[282]=25'd375;
            NN[283]=-25'd1093;
            NN[284]=-25'd2967;
            NN[285]=-25'd3697;
            NN[286]=-25'd6286;
            NN[287]=-25'd5696;
            NN[288]=-25'd4234;
            NN[289]=25'd261;
            NN[290]=-25'd2910;
            NN[291]=25'd2323;
            NN[292]=25'd5066;
            NN[293]=25'd6337;
            NN[294]=-25'd2182;
            NN[295]=-25'd11148;
            NN[296]=-25'd5394;
            NN[297]=25'd10984;
            NN[298]=25'd17590;
            NN[299]=25'd14096;
            NN[300]=25'd14254;
            NN[301]=25'd10359;
            NN[302]=25'd19941;
            NN[303]=25'd29028;
            NN[304]=25'd11879;
            NN[305]=-25'd7051;
            NN[306]=-25'd2986;
            NN[307]=-25'd44;
            NN[308]=-25'd1;
            NN[309]=25'd109;
            NN[310]=-25'd229;
            NN[311]=-25'd1435;
            NN[312]=-25'd5731;
            NN[313]=-25'd4769;
            NN[314]=-25'd2420;
            NN[315]=-25'd992;
            NN[316]=-25'd1707;
            NN[317]=-25'd3013;
            NN[318]=-25'd1147;
            NN[319]=25'd1014;
            NN[320]=-25'd1538;
            NN[321]=-25'd5151;
            NN[322]=-25'd27090;
            NN[323]=-25'd41886;
            NN[324]=-25'd37709;
            NN[325]=-25'd12232;
            NN[326]=-25'd981;
            NN[327]=25'd9183;
            NN[328]=25'd12680;
            NN[329]=25'd16448;
            NN[330]=25'd25517;
            NN[331]=25'd30450;
            NN[332]=25'd17010;
            NN[333]=-25'd2763;
            NN[334]=-25'd1515;
            NN[335]=-25'd36;
            NN[336]=-25'd1;
            NN[337]=-25'd2;
            NN[338]=-25'd205;
            NN[339]=-25'd1760;
            NN[340]=-25'd5652;
            NN[341]=-25'd1753;
            NN[342]=25'd6034;
            NN[343]=25'd4348;
            NN[344]=25'd217;
            NN[345]=25'd993;
            NN[346]=25'd5112;
            NN[347]=25'd4921;
            NN[348]=25'd3306;
            NN[349]=-25'd14115;
            NN[350]=-25'd44406;
            NN[351]=-25'd57495;
            NN[352]=-25'd50798;
            NN[353]=-25'd23534;
            NN[354]=-25'd7285;
            NN[355]=25'd1714;
            NN[356]=25'd1481;
            NN[357]=25'd11526;
            NN[358]=25'd30437;
            NN[359]=25'd32935;
            NN[360]=25'd21851;
            NN[361]=25'd692;
            NN[362]=-25'd471;
            NN[363]=-25'd9;
            NN[364]=25'd0;
            NN[365]=25'd39;
            NN[366]=-25'd111;
            NN[367]=-25'd1346;
            NN[368]=-25'd3881;
            NN[369]=25'd815;
            NN[370]=25'd12192;
            NN[371]=25'd14937;
            NN[372]=25'd8334;
            NN[373]=25'd9474;
            NN[374]=25'd13040;
            NN[375]=25'd9450;
            NN[376]=25'd1551;
            NN[377]=-25'd30513;
            NN[378]=-25'd52048;
            NN[379]=-25'd60154;
            NN[380]=-25'd52241;
            NN[381]=-25'd27943;
            NN[382]=-25'd9933;
            NN[383]=-25'd9211;
            NN[384]=-25'd11027;
            NN[385]=25'd8779;
            NN[386]=25'd28703;
            NN[387]=25'd31243;
            NN[388]=25'd19407;
            NN[389]=25'd1644;
            NN[390]=-25'd200;
            NN[391]=-25'd51;
        end
        1:begin
            NN[0]=-25'd9;
            NN[1]=-25'd9;
            NN[2]=-25'd59;
            NN[3]=-25'd2141;
            NN[4]=-25'd3656;
            NN[5]=25'd8592;
            NN[6]=25'd16013;
            NN[7]=25'd21889;
            NN[8]=25'd17307;
            NN[9]=25'd17018;
            NN[10]=25'd14987;
            NN[11]=25'd10967;
            NN[12]=-25'd5213;
            NN[13]=-25'd35369;
            NN[14]=-25'd55183;
            NN[15]=-25'd58193;
            NN[16]=-25'd51778;
            NN[17]=-25'd23642;
            NN[18]=-25'd9843;
            NN[19]=-25'd10613;
            NN[20]=-25'd3834;
            NN[21]=25'd12676;
            NN[22]=25'd22432;
            NN[23]=25'd26826;
            NN[24]=25'd17985;
            NN[25]=25'd616;
            NN[26]=-25'd244;
            NN[27]=-25'd10;
            NN[28]=-25'd3;
            NN[29]=-25'd20;
            NN[30]=-25'd87;
            NN[31]=-25'd2469;
            NN[32]=-25'd158;
            NN[33]=25'd15992;
            NN[34]=25'd17525;
            NN[35]=25'd22540;
            NN[36]=25'd19878;
            NN[37]=25'd21758;
            NN[38]=25'd20390;
            NN[39]=25'd2816;
            NN[40]=-25'd19321;
            NN[41]=-25'd48900;
            NN[42]=-25'd61267;
            NN[43]=-25'd56315;
            NN[44]=-25'd40608;
            NN[45]=-25'd19688;
            NN[46]=-25'd6318;
            NN[47]=-25'd3149;
            NN[48]=25'd5616;
            NN[49]=25'd11498;
            NN[50]=25'd20085;
            NN[51]=25'd22985;
            NN[52]=25'd13322;
            NN[53]=-25'd382;
            NN[54]=-25'd314;
            NN[55]=-25'd43;
            NN[56]=25'd0;
            NN[57]=-25'd10;
            NN[58]=-25'd139;
            NN[59]=-25'd2506;
            NN[60]=25'd1605;
            NN[61]=25'd19995;
            NN[62]=25'd23770;
            NN[63]=25'd18324;
            NN[64]=25'd20380;
            NN[65]=25'd21311;
            NN[66]=25'd21427;
            NN[67]=25'd918;
            NN[68]=-25'd28674;
            NN[69]=-25'd54102;
            NN[70]=-25'd57021;
            NN[71]=-25'd46597;
            NN[72]=-25'd27605;
            NN[73]=-25'd7462;
            NN[74]=25'd185;
            NN[75]=25'd3321;
            NN[76]=25'd8922;
            NN[77]=25'd12856;
            NN[78]=25'd16256;
            NN[79]=25'd15511;
            NN[80]=25'd4580;
            NN[81]=-25'd2250;
            NN[82]=-25'd827;
            NN[83]=-25'd25;
            NN[84]=25'd0;
            NN[85]=-25'd4;
            NN[86]=-25'd282;
            NN[87]=-25'd3321;
            NN[88]=25'd876;
            NN[89]=25'd17226;
            NN[90]=25'd21495;
            NN[91]=25'd16695;
            NN[92]=25'd14932;
            NN[93]=25'd21274;
            NN[94]=25'd24027;
            NN[95]=-25'd1481;
            NN[96]=-25'd26692;
            NN[97]=-25'd50360;
            NN[98]=-25'd51160;
            NN[99]=-25'd33496;
            NN[100]=-25'd10862;
            NN[101]=25'd2536;
            NN[102]=25'd455;
            NN[103]=25'd2343;
            NN[104]=25'd5138;
            NN[105]=25'd6574;
            NN[106]=25'd14916;
            NN[107]=25'd7801;
            NN[108]=-25'd19;
            NN[109]=-25'd1719;
            NN[110]=-25'd534;
            NN[111]=25'd335;
            NN[112]=-25'd3;
            NN[113]=25'd0;
            NN[114]=-25'd248;
            NN[115]=-25'd5490;
            NN[116]=-25'd1273;
            NN[117]=25'd11848;
            NN[118]=25'd15654;
            NN[119]=25'd14381;
            NN[120]=25'd16739;
            NN[121]=25'd21714;
            NN[122]=25'd24412;
            NN[123]=25'd3110;
            NN[124]=-25'd22744;
            NN[125]=-25'd39564;
            NN[126]=-25'd37024;
            NN[127]=-25'd19486;
            NN[128]=-25'd5049;
            NN[129]=25'd338;
            NN[130]=-25'd2386;
            NN[131]=-25'd604;
            NN[132]=-25'd2654;
            NN[133]=25'd5022;
            NN[134]=25'd11339;
            NN[135]=25'd3590;
            NN[136]=-25'd2185;
            NN[137]=-25'd1623;
            NN[138]=-25'd411;
            NN[139]=-25'd202;
            NN[140]=25'd0;
            NN[141]=25'd149;
            NN[142]=-25'd148;
            NN[143]=-25'd4833;
            NN[144]=-25'd2359;
            NN[145]=25'd8365;
            NN[146]=25'd16191;
            NN[147]=25'd14776;
            NN[148]=25'd14885;
            NN[149]=25'd19696;
            NN[150]=25'd27071;
            NN[151]=25'd18856;
            NN[152]=25'd3467;
            NN[153]=-25'd12375;
            NN[154]=-25'd14712;
            NN[155]=-25'd8948;
            NN[156]=-25'd5394;
            NN[157]=-25'd905;
            NN[158]=-25'd3499;
            NN[159]=-25'd6200;
            NN[160]=-25'd1919;
            NN[161]=25'd4318;
            NN[162]=25'd6281;
            NN[163]=-25'd1534;
            NN[164]=-25'd2248;
            NN[165]=-25'd1523;
            NN[166]=-25'd322;
            NN[167]=-25'd56;
            NN[168]=25'd0;
            NN[169]=25'd378;
            NN[170]=-25'd39;
            NN[171]=-25'd3822;
            NN[172]=-25'd2139;
            NN[173]=25'd10821;
            NN[174]=25'd14836;
            NN[175]=25'd13100;
            NN[176]=25'd9762;
            NN[177]=25'd16605;
            NN[178]=25'd28845;
            NN[179]=25'd30293;
            NN[180]=25'd19993;
            NN[181]=25'd6734;
            NN[182]=-25'd290;
            NN[183]=-25'd438;
            NN[184]=-25'd4759;
            NN[185]=-25'd3300;
            NN[186]=-25'd8044;
            NN[187]=-25'd9202;
            NN[188]=-25'd3856;
            NN[189]=25'd1532;
            NN[190]=-25'd534;
            NN[191]=-25'd3833;
            NN[192]=-25'd2388;
            NN[193]=-25'd908;
            NN[194]=-25'd84;
            NN[195]=25'd0;
            NN[196]=25'd0;
            NN[197]=-25'd2;
            NN[198]=-25'd170;
            NN[199]=-25'd2653;
            NN[200]=-25'd4134;
            NN[201]=25'd6480;
            NN[202]=25'd11852;
            NN[203]=25'd12225;
            NN[204]=25'd5261;
            NN[205]=25'd10616;
            NN[206]=25'd21772;
            NN[207]=25'd28155;
            NN[208]=25'd18993;
            NN[209]=25'd7134;
            NN[210]=25'd1413;
            NN[211]=-25'd1003;
            NN[212]=-25'd520;
            NN[213]=-25'd4914;
            NN[214]=-25'd8492;
            NN[215]=-25'd10831;
            NN[216]=-25'd5604;
            NN[217]=-25'd4053;
            NN[218]=-25'd3871;
            NN[219]=-25'd2443;
            NN[220]=-25'd1519;
            NN[221]=-25'd322;
            NN[222]=25'd130;
            NN[223]=25'd0;
            NN[224]=25'd0;
            NN[225]=25'd0;
            NN[226]=-25'd102;
            NN[227]=-25'd2058;
            NN[228]=-25'd6772;
            NN[229]=-25'd443;
            NN[230]=25'd7170;
            NN[231]=25'd9849;
            NN[232]=25'd13992;
            NN[233]=25'd14403;
            NN[234]=25'd18094;
            NN[235]=25'd24357;
            NN[236]=25'd21006;
            NN[237]=25'd23332;
            NN[238]=25'd13587;
            NN[239]=25'd10386;
            NN[240]=25'd6793;
            NN[241]=25'd429;
            NN[242]=-25'd8157;
            NN[243]=-25'd11182;
            NN[244]=-25'd12248;
            NN[245]=-25'd8350;
            NN[246]=-25'd3197;
            NN[247]=-25'd796;
            NN[248]=-25'd604;
            NN[249]=-25'd88;
            NN[250]=25'd16;
            NN[251]=25'd0;
            NN[252]=25'd0;
            NN[253]=25'd0;
            NN[254]=-25'd18;
            NN[255]=-25'd844;
            NN[256]=-25'd4249;
            NN[257]=-25'd4884;
            NN[258]=-25'd392;
            NN[259]=25'd5079;
            NN[260]=25'd10037;
            NN[261]=25'd14806;
            NN[262]=25'd18958;
            NN[263]=25'd24893;
            NN[264]=25'd26702;
            NN[265]=25'd25992;
            NN[266]=25'd20918;
            NN[267]=25'd12962;
            NN[268]=25'd2483;
            NN[269]=-25'd3946;
            NN[270]=-25'd16192;
            NN[271]=-25'd16823;
            NN[272]=-25'd13330;
            NN[273]=-25'd7033;
            NN[274]=-25'd3097;
            NN[275]=-25'd1180;
            NN[276]=-25'd478;
            NN[277]=-25'd28;
            NN[278]=25'd0;
            NN[279]=25'd0;
            NN[280]=25'd0;
            NN[281]=25'd0;
            NN[282]=-25'd73;
            NN[283]=-25'd123;
            NN[284]=-25'd743;
            NN[285]=-25'd2414;
            NN[286]=-25'd3512;
            NN[287]=-25'd6400;
            NN[288]=-25'd5227;
            NN[289]=-25'd4377;
            NN[290]=-25'd3196;
            NN[291]=-25'd1709;
            NN[292]=25'd5280;
            NN[293]=25'd5364;
            NN[294]=25'd1224;
            NN[295]=-25'd4612;
            NN[296]=-25'd8558;
            NN[297]=-25'd11856;
            NN[298]=-25'd13200;
            NN[299]=-25'd11039;
            NN[300]=-25'd8767;
            NN[301]=-25'd5857;
            NN[302]=-25'd2570;
            NN[303]=-25'd875;
            NN[304]=-25'd101;
            NN[305]=-25'd9;
            NN[306]=25'd0;
            NN[307]=25'd0;
            NN[308]=25'd0;
            NN[309]=25'd0;
            NN[310]=25'd0;
            NN[311]=-25'd4;
            NN[312]=-25'd129;
            NN[313]=-25'd549;
            NN[314]=-25'd2182;
            NN[315]=-25'd4510;
            NN[316]=-25'd7633;
            NN[317]=-25'd11613;
            NN[318]=-25'd14294;
            NN[319]=-25'd14879;
            NN[320]=-25'd17203;
            NN[321]=-25'd16652;
            NN[322]=-25'd15143;
            NN[323]=-25'd13234;
            NN[324]=-25'd10617;
            NN[325]=-25'd9874;
            NN[326]=-25'd7770;
            NN[327]=-25'd5518;
            NN[328]=-25'd4644;
            NN[329]=-25'd3153;
            NN[330]=-25'd1267;
            NN[331]=-25'd305;
            NN[332]=-25'd51;
            NN[333]=25'd0;
            NN[334]=25'd0;
            NN[335]=25'd0;
            NN[336]=25'd0;
            NN[337]=25'd0;
            NN[338]=25'd0;
            NN[339]=25'd0;
            NN[340]=-25'd15;
            NN[341]=-25'd168;
            NN[342]=-25'd560;
            NN[343]=-25'd1386;
            NN[344]=-25'd2145;
            NN[345]=-25'd3627;
            NN[346]=-25'd3195;
            NN[347]=-25'd2874;
            NN[348]=-25'd2518;
            NN[349]=-25'd3703;
            NN[350]=-25'd4460;
            NN[351]=-25'd3638;
            NN[352]=-25'd3086;
            NN[353]=-25'd2820;
            NN[354]=-25'd1989;
            NN[355]=-25'd671;
            NN[356]=-25'd1037;
            NN[357]=-25'd1047;
            NN[358]=-25'd628;
            NN[359]=-25'd48;
            NN[360]=25'd0;
            NN[361]=25'd0;
            NN[362]=25'd0;
            NN[363]=25'd0;
            NN[364]=25'd0;
            NN[365]=25'd0;
            NN[366]=25'd0;
            NN[367]=25'd0;
            NN[368]=25'd0;
            NN[369]=-25'd1;
            NN[370]=-25'd4;
            NN[371]=-25'd25;
            NN[372]=-25'd77;
            NN[373]=-25'd141;
            NN[374]=-25'd89;
            NN[375]=-25'd155;
            NN[376]=-25'd246;
            NN[377]=-25'd325;
            NN[378]=-25'd585;
            NN[379]=-25'd667;
            NN[380]=-25'd523;
            NN[381]=-25'd341;
            NN[382]=-25'd257;
            NN[383]=-25'd119;
            NN[384]=-25'd199;
            NN[385]=-25'd261;
            NN[386]=-25'd682;
            NN[387]=-25'd157;
            NN[388]=25'd0;
            NN[389]=25'd0;
            NN[390]=25'd0;
            NN[391]=25'd0;
        end
        2:begin
            NN[0]=25'd0;
            NN[1]=25'd0;
            NN[2]=25'd0;
            NN[3]=25'd0;
            NN[4]=25'd0;
            NN[5]=25'd0;
            NN[6]=25'd0;
            NN[7]=25'd0;
            NN[8]=25'd0;
            NN[9]=25'd0;
            NN[10]=25'd0;
            NN[11]=25'd0;
            NN[12]=25'd0;
            NN[13]=25'd0;
            NN[14]=25'd0;
            NN[15]=25'd0;
            NN[16]=25'd0;
            NN[17]=25'd0;
            NN[18]=25'd0;
            NN[19]=25'd0;
            NN[20]=25'd0;
            NN[21]=25'd0;
            NN[22]=25'd0;
            NN[23]=25'd0;
            NN[24]=25'd0;
            NN[25]=25'd0;
            NN[26]=25'd0;
            NN[27]=25'd0;
            NN[28]=25'd0;
            NN[29]=25'd0;
            NN[30]=25'd0;
            NN[31]=25'd0;
            NN[32]=25'd0;
            NN[33]=25'd0;
            NN[34]=25'd0;
            NN[35]=-25'd1;
            NN[36]=-25'd65;
            NN[37]=-25'd82;
            NN[38]=-25'd127;
            NN[39]=-25'd56;
            NN[40]=-25'd44;
            NN[41]=-25'd23;
            NN[42]=25'd385;
            NN[43]=25'd649;
            NN[44]=-25'd186;
            NN[45]=-25'd105;
            NN[46]=-25'd10;
            NN[47]=-25'd10;
            NN[48]=-25'd10;
            NN[49]=-25'd8;
            NN[50]=25'd0;
            NN[51]=25'd0;
            NN[52]=25'd0;
            NN[53]=25'd0;
            NN[54]=25'd0;
            NN[55]=25'd0;
            NN[56]=25'd0;
            NN[57]=25'd0;
            NN[58]=25'd0;
            NN[59]=25'd0;
            NN[60]=25'd0;
            NN[61]=25'd0;
            NN[62]=-25'd1;
            NN[63]=-25'd58;
            NN[64]=-25'd556;
            NN[65]=-25'd1154;
            NN[66]=-25'd1161;
            NN[67]=-25'd1316;
            NN[68]=-25'd321;
            NN[69]=25'd2198;
            NN[70]=25'd2952;
            NN[71]=25'd4964;
            NN[72]=25'd2764;
            NN[73]=25'd166;
            NN[74]=-25'd509;
            NN[75]=25'd16;
            NN[76]=-25'd455;
            NN[77]=-25'd498;
            NN[78]=-25'd374;
            NN[79]=-25'd124;
            NN[80]=-25'd34;
            NN[81]=-25'd5;
            NN[82]=25'd0;
            NN[83]=25'd0;
            NN[84]=25'd0;
            NN[85]=25'd0;
            NN[86]=25'd8;
            NN[87]=25'd2;
            NN[88]=-25'd2;
            NN[89]=-25'd46;
            NN[90]=-25'd99;
            NN[91]=-25'd625;
            NN[92]=-25'd2184;
            NN[93]=-25'd3500;
            NN[94]=-25'd5180;
            NN[95]=-25'd7479;
            NN[96]=-25'd4695;
            NN[97]=-25'd1378;
            NN[98]=25'd13;
            NN[99]=25'd2677;
            NN[100]=25'd1424;
            NN[101]=-25'd2720;
            NN[102]=-25'd5444;
            NN[103]=-25'd4565;
            NN[104]=-25'd4394;
            NN[105]=-25'd3587;
            NN[106]=-25'd2393;
            NN[107]=-25'd1439;
            NN[108]=-25'd974;
            NN[109]=-25'd258;
            NN[110]=-25'd348;
            NN[111]=25'd0;
            NN[112]=25'd0;
            NN[113]=25'd0;
            NN[114]=25'd28;
            NN[115]=-25'd1;
            NN[116]=25'd68;
            NN[117]=25'd581;
            NN[118]=-25'd243;
            NN[119]=-25'd2528;
            NN[120]=-25'd4813;
            NN[121]=-25'd6772;
            NN[122]=-25'd6438;
            NN[123]=-25'd6734;
            NN[124]=25'd210;
            NN[125]=25'd11429;
            NN[126]=25'd16353;
            NN[127]=25'd12278;
            NN[128]=25'd6719;
            NN[129]=25'd1799;
            NN[130]=-25'd561;
            NN[131]=25'd6854;
            NN[132]=25'd9875;
            NN[133]=25'd9002;
            NN[134]=25'd5174;
            NN[135]=25'd1594;
            NN[136]=-25'd3059;
            NN[137]=-25'd1810;
            NN[138]=-25'd204;
            NN[139]=-25'd79;
            NN[140]=25'd0;
            NN[141]=25'd0;
            NN[142]=25'd2;
            NN[143]=25'd120;
            NN[144]=25'd148;
            NN[145]=25'd710;
            NN[146]=-25'd1982;
            NN[147]=-25'd6801;
            NN[148]=-25'd12978;
            NN[149]=-25'd14541;
            NN[150]=-25'd10549;
            NN[151]=-25'd7361;
            NN[152]=25'd371;
            NN[153]=25'd8674;
            NN[154]=25'd11922;
            NN[155]=25'd10748;
            NN[156]=-25'd2556;
            NN[157]=-25'd7156;
            NN[158]=-25'd847;
            NN[159]=25'd6981;
            NN[160]=25'd14088;
            NN[161]=25'd17994;
            NN[162]=25'd15333;
            NN[163]=25'd7393;
            NN[164]=25'd851;
            NN[165]=-25'd2693;
            NN[166]=-25'd343;
            NN[167]=-25'd90;
            NN[168]=25'd0;
            NN[169]=25'd0;
            NN[170]=-25'd263;
            NN[171]=25'd32;
            NN[172]=25'd13;
            NN[173]=-25'd2174;
            NN[174]=-25'd5657;
            NN[175]=-25'd11627;
            NN[176]=-25'd18768;
            NN[177]=-25'd23304;
            NN[178]=-25'd16998;
            NN[179]=-25'd10765;
            NN[180]=-25'd8355;
            NN[181]=-25'd7931;
            NN[182]=-25'd8932;
            NN[183]=-25'd14408;
            NN[184]=-25'd17345;
            NN[185]=-25'd17757;
            NN[186]=-25'd8172;
            NN[187]=-25'd1813;
            NN[188]=25'd9190;
            NN[189]=25'd10136;
            NN[190]=25'd8185;
            NN[191]=25'd3222;
            NN[192]=-25'd1645;
            NN[193]=-25'd3142;
            NN[194]=-25'd298;
            NN[195]=-25'd14;
            NN[196]=25'd0;
            NN[197]=-25'd8;
            NN[198]=-25'd244;
            NN[199]=-25'd357;
            NN[200]=-25'd606;
            NN[201]=-25'd4219;
            NN[202]=-25'd9398;
            NN[203]=-25'd14053;
            NN[204]=-25'd23910;
            NN[205]=-25'd25963;
            NN[206]=-25'd23151;
            NN[207]=-25'd18996;
            NN[208]=-25'd12273;
            NN[209]=-25'd12549;
            NN[210]=-25'd13605;
            NN[211]=-25'd22055;
            NN[212]=-25'd20764;
            NN[213]=-25'd16442;
            NN[214]=-25'd12464;
            NN[215]=-25'd2374;
            NN[216]=25'd3382;
            NN[217]=-25'd149;
            NN[218]=-25'd1305;
            NN[219]=-25'd5922;
            NN[220]=-25'd9979;
            NN[221]=-25'd5505;
            NN[222]=-25'd443;
            NN[223]=-25'd122;
            NN[224]=25'd0;
            NN[225]=-25'd10;
            NN[226]=-25'd123;
            NN[227]=-25'd261;
            NN[228]=-25'd852;
            NN[229]=-25'd4020;
            NN[230]=-25'd9221;
            NN[231]=-25'd13159;
            NN[232]=-25'd22654;
            NN[233]=-25'd27673;
            NN[234]=-25'd25039;
            NN[235]=-25'd19046;
            NN[236]=-25'd10051;
            NN[237]=-25'd3905;
            NN[238]=-25'd1879;
            NN[239]=25'd762;
            NN[240]=-25'd9589;
            NN[241]=25'd306;
            NN[242]=-25'd5767;
            NN[243]=-25'd5260;
            NN[244]=-25'd8510;
            NN[245]=-25'd13625;
            NN[246]=-25'd16715;
            NN[247]=-25'd18825;
            NN[248]=-25'd16092;
            NN[249]=-25'd7420;
            NN[250]=-25'd820;
            NN[251]=-25'd95;
            NN[252]=25'd0;
            NN[253]=-25'd1;
            NN[254]=-25'd59;
            NN[255]=-25'd272;
            NN[256]=-25'd1466;
            NN[257]=-25'd6024;
            NN[258]=-25'd8679;
            NN[259]=-25'd11145;
            NN[260]=-25'd17747;
            NN[261]=-25'd22952;
            NN[262]=-25'd19430;
            NN[263]=-25'd12084;
            NN[264]=-25'd6508;
            NN[265]=25'd5857;
            NN[266]=25'd20591;
            NN[267]=25'd29201;
            NN[268]=25'd11533;
            NN[269]=25'd1773;
            NN[270]=-25'd7257;
            NN[271]=-25'd15318;
            NN[272]=-25'd20537;
            NN[273]=-25'd23254;
            NN[274]=-25'd24324;
            NN[275]=-25'd21727;
            NN[276]=-25'd14088;
            NN[277]=-25'd5776;
            NN[278]=-25'd750;
            NN[279]=-25'd71;
            NN[280]=25'd0;
            NN[281]=-25'd1;
            NN[282]=-25'd30;
            NN[283]=-25'd786;
            NN[284]=-25'd1708;
            NN[285]=-25'd5960;
            NN[286]=-25'd10195;
            NN[287]=-25'd11075;
            NN[288]=-25'd13732;
            NN[289]=-25'd18180;
            NN[290]=-25'd13902;
            NN[291]=-25'd8302;
            NN[292]=-25'd2318;
            NN[293]=25'd15876;
            NN[294]=25'd44001;
            NN[295]=25'd50116;
            NN[296]=25'd19651;
            NN[297]=25'd638;
            NN[298]=-25'd13768;
            NN[299]=-25'd17913;
            NN[300]=-25'd23875;
            NN[301]=-25'd21805;
            NN[302]=-25'd19593;
            NN[303]=-25'd15926;
            NN[304]=-25'd10639;
            NN[305]=-25'd3552;
            NN[306]=-25'd674;
            NN[307]=25'd35;
            NN[308]=25'd0;
            NN[309]=25'd5;
            NN[310]=-25'd11;
            NN[311]=-25'd552;
            NN[312]=-25'd889;
            NN[313]=-25'd3679;
            NN[314]=-25'd8564;
            NN[315]=-25'd10599;
            NN[316]=-25'd12364;
            NN[317]=-25'd16731;
            NN[318]=-25'd16562;
            NN[319]=-25'd16448;
            NN[320]=-25'd6495;
            NN[321]=25'd19597;
            NN[322]=25'd58922;
            NN[323]=25'd56756;
            NN[324]=25'd16682;
            NN[325]=-25'd4697;
            NN[326]=-25'd10675;
            NN[327]=-25'd16621;
            NN[328]=-25'd16817;
            NN[329]=-25'd13869;
            NN[330]=-25'd10239;
            NN[331]=-25'd7506;
            NN[332]=-25'd5255;
            NN[333]=-25'd2297;
            NN[334]=-25'd433;
            NN[335]=25'd54;
            NN[336]=25'd0;
            NN[337]=-25'd3;
            NN[338]=-25'd43;
            NN[339]=-25'd116;
            NN[340]=-25'd127;
            NN[341]=-25'd2732;
            NN[342]=-25'd5076;
            NN[343]=-25'd7121;
            NN[344]=-25'd10670;
            NN[345]=-25'd14302;
            NN[346]=-25'd24219;
            NN[347]=-25'd30651;
            NN[348]=-25'd9589;
            NN[349]=25'd23035;
            NN[350]=25'd70925;
            NN[351]=25'd49349;
            NN[352]=25'd10261;
            NN[353]=25'd287;
            NN[354]=-25'd10053;
            NN[355]=-25'd15654;
            NN[356]=-25'd12179;
            NN[357]=-25'd7437;
            NN[358]=-25'd5431;
            NN[359]=-25'd3284;
            NN[360]=-25'd2287;
            NN[361]=-25'd859;
            NN[362]=-25'd372;
            NN[363]=25'd22;
            NN[364]=25'd2;
            NN[365]=25'd0;
            NN[366]=-25'd14;
            NN[367]=25'd48;
            NN[368]=25'd6;
            NN[369]=-25'd2355;
            NN[370]=-25'd4653;
            NN[371]=-25'd7017;
            NN[372]=-25'd7601;
            NN[373]=-25'd17026;
            NN[374]=-25'd35258;
            NN[375]=-25'd40803;
            NN[376]=-25'd16044;
            NN[377]=25'd30874;
            NN[378]=25'd63218;
            NN[379]=25'd40862;
            NN[380]=25'd9624;
            NN[381]=-25'd3098;
            NN[382]=-25'd19335;
            NN[383]=-25'd16869;
            NN[384]=-25'd11174;
            NN[385]=-25'd7341;
            NN[386]=-25'd5802;
            NN[387]=-25'd4650;
            NN[388]=-25'd3372;
            NN[389]=-25'd1408;
            NN[390]=-25'd586;
            NN[391]=-25'd24;
        end
        3:begin
            NN[0]=25'd0;
            NN[1]=-25'd1;
            NN[2]=25'd6;
            NN[3]=25'd116;
            NN[4]=25'd188;
            NN[5]=-25'd2761;
            NN[6]=-25'd5292;
            NN[7]=-25'd8142;
            NN[8]=-25'd9395;
            NN[9]=-25'd20579;
            NN[10]=-25'd38975;
            NN[11]=-25'd41515;
            NN[12]=-25'd7241;
            NN[13]=25'd34985;
            NN[14]=25'd55135;
            NN[15]=25'd35235;
            NN[16]=25'd3277;
            NN[17]=-25'd22723;
            NN[18]=-25'd29920;
            NN[19]=-25'd21850;
            NN[20]=-25'd14273;
            NN[21]=-25'd9286;
            NN[22]=-25'd6604;
            NN[23]=-25'd4860;
            NN[24]=-25'd2577;
            NN[25]=-25'd1258;
            NN[26]=-25'd266;
            NN[27]=-25'd23;
            NN[28]=25'd0;
            NN[29]=-25'd2;
            NN[30]=25'd78;
            NN[31]=25'd79;
            NN[32]=-25'd370;
            NN[33]=-25'd4078;
            NN[34]=-25'd8215;
            NN[35]=-25'd9539;
            NN[36]=-25'd11764;
            NN[37]=-25'd22684;
            NN[38]=-25'd32969;
            NN[39]=-25'd22180;
            NN[40]=25'd3484;
            NN[41]=25'd38352;
            NN[42]=25'd54585;
            NN[43]=25'd19940;
            NN[44]=-25'd8580;
            NN[45]=-25'd34654;
            NN[46]=-25'd31411;
            NN[47]=-25'd23866;
            NN[48]=-25'd16396;
            NN[49]=-25'd10780;
            NN[50]=-25'd7819;
            NN[51]=-25'd5306;
            NN[52]=-25'd3157;
            NN[53]=-25'd1348;
            NN[54]=-25'd500;
            NN[55]=-25'd102;
            NN[56]=25'd0;
            NN[57]=25'd1;
            NN[58]=25'd133;
            NN[59]=-25'd134;
            NN[60]=-25'd836;
            NN[61]=-25'd5781;
            NN[62]=-25'd13214;
            NN[63]=-25'd16397;
            NN[64]=-25'd18166;
            NN[65]=-25'd17967;
            NN[66]=-25'd13647;
            NN[67]=-25'd11047;
            NN[68]=-25'd1926;
            NN[69]=25'd36930;
            NN[70]=25'd49987;
            NN[71]=25'd4838;
            NN[72]=-25'd20647;
            NN[73]=-25'd40010;
            NN[74]=-25'd33034;
            NN[75]=-25'd23456;
            NN[76]=-25'd15763;
            NN[77]=-25'd10897;
            NN[78]=-25'd8476;
            NN[79]=-25'd6463;
            NN[80]=-25'd4093;
            NN[81]=-25'd2485;
            NN[82]=-25'd921;
            NN[83]=-25'd20;
            NN[84]=25'd0;
            NN[85]=25'd27;
            NN[86]=-25'd23;
            NN[87]=-25'd341;
            NN[88]=-25'd1700;
            NN[89]=-25'd10172;
            NN[90]=-25'd19849;
            NN[91]=-25'd22534;
            NN[92]=-25'd19746;
            NN[93]=-25'd12001;
            NN[94]=25'd521;
            NN[95]=-25'd4982;
            NN[96]=25'd7976;
            NN[97]=25'd36536;
            NN[98]=25'd34113;
            NN[99]=-25'd2433;
            NN[100]=-25'd25826;
            NN[101]=-25'd34243;
            NN[102]=-25'd26587;
            NN[103]=-25'd18062;
            NN[104]=-25'd12138;
            NN[105]=-25'd9004;
            NN[106]=-25'd6765;
            NN[107]=-25'd5981;
            NN[108]=-25'd4042;
            NN[109]=-25'd3015;
            NN[110]=-25'd582;
            NN[111]=-25'd20;
            NN[112]=-25'd3;
            NN[113]=25'd4;
            NN[114]=-25'd49;
            NN[115]=-25'd453;
            NN[116]=-25'd3170;
            NN[117]=-25'd12998;
            NN[118]=-25'd24719;
            NN[119]=-25'd24553;
            NN[120]=-25'd12512;
            NN[121]=-25'd2087;
            NN[122]=-25'd2986;
            NN[123]=-25'd1865;
            NN[124]=25'd10253;
            NN[125]=25'd23344;
            NN[126]=25'd17428;
            NN[127]=-25'd9088;
            NN[128]=-25'd21851;
            NN[129]=-25'd17851;
            NN[130]=-25'd13218;
            NN[131]=-25'd9454;
            NN[132]=-25'd5884;
            NN[133]=-25'd5566;
            NN[134]=-25'd6353;
            NN[135]=-25'd5681;
            NN[136]=-25'd2497;
            NN[137]=-25'd419;
            NN[138]=25'd48;
            NN[139]=-25'd4;
            NN[140]=25'd2;
            NN[141]=25'd12;
            NN[142]=-25'd50;
            NN[143]=-25'd600;
            NN[144]=-25'd4274;
            NN[145]=-25'd15628;
            NN[146]=-25'd18555;
            NN[147]=-25'd14065;
            NN[148]=-25'd6302;
            NN[149]=25'd1222;
            NN[150]=-25'd4117;
            NN[151]=25'd675;
            NN[152]=25'd1748;
            NN[153]=25'd14791;
            NN[154]=25'd2936;
            NN[155]=-25'd5270;
            NN[156]=-25'd2593;
            NN[157]=-25'd3303;
            NN[158]=-25'd1770;
            NN[159]=-25'd210;
            NN[160]=-25'd2716;
            NN[161]=-25'd3726;
            NN[162]=-25'd5139;
            NN[163]=-25'd3576;
            NN[164]=-25'd500;
            NN[165]=25'd914;
            NN[166]=25'd41;
            NN[167]=25'd0;
            NN[168]=25'd0;
            NN[169]=-25'd2;
            NN[170]=-25'd271;
            NN[171]=-25'd1007;
            NN[172]=-25'd2874;
            NN[173]=-25'd9694;
            NN[174]=-25'd5574;
            NN[175]=-25'd1449;
            NN[176]=25'd6364;
            NN[177]=25'd6021;
            NN[178]=25'd5596;
            NN[179]=25'd5026;
            NN[180]=-25'd294;
            NN[181]=-25'd145;
            NN[182]=-25'd458;
            NN[183]=-25'd4116;
            NN[184]=25'd6994;
            NN[185]=25'd12314;
            NN[186]=25'd10395;
            NN[187]=25'd5400;
            NN[188]=25'd800;
            NN[189]=-25'd2895;
            NN[190]=-25'd4583;
            NN[191]=-25'd4134;
            NN[192]=-25'd2445;
            NN[193]=-25'd249;
            NN[194]=25'd84;
            NN[195]=25'd9;
            NN[196]=25'd2;
            NN[197]=25'd0;
            NN[198]=-25'd492;
            NN[199]=-25'd581;
            NN[200]=25'd1331;
            NN[201]=25'd8877;
            NN[202]=25'd10135;
            NN[203]=25'd9086;
            NN[204]=25'd11813;
            NN[205]=25'd6682;
            NN[206]=25'd7434;
            NN[207]=-25'd7708;
            NN[208]=-25'd13555;
            NN[209]=-25'd12675;
            NN[210]=-25'd3636;
            NN[211]=25'd714;
            NN[212]=25'd6205;
            NN[213]=25'd11229;
            NN[214]=25'd12312;
            NN[215]=25'd5533;
            NN[216]=25'd1816;
            NN[217]=-25'd1160;
            NN[218]=-25'd6965;
            NN[219]=-25'd5158;
            NN[220]=-25'd1379;
            NN[221]=-25'd379;
            NN[222]=-25'd109;
            NN[223]=25'd0;
            NN[224]=25'd1;
            NN[225]=25'd0;
            NN[226]=-25'd497;
            NN[227]=-25'd466;
            NN[228]=25'd3640;
            NN[229]=25'd19811;
            NN[230]=25'd18903;
            NN[231]=25'd13865;
            NN[232]=25'd9546;
            NN[233]=25'd6831;
            NN[234]=-25'd3129;
            NN[235]=-25'd21223;
            NN[236]=-25'd28913;
            NN[237]=-25'd23989;
            NN[238]=-25'd9586;
            NN[239]=25'd2122;
            NN[240]=25'd9089;
            NN[241]=25'd16191;
            NN[242]=25'd12091;
            NN[243]=25'd3589;
            NN[244]=-25'd465;
            NN[245]=-25'd4533;
            NN[246]=-25'd5758;
            NN[247]=-25'd3119;
            NN[248]=-25'd908;
            NN[249]=-25'd143;
            NN[250]=25'd142;
            NN[251]=25'd0;
            NN[252]=25'd0;
            NN[253]=25'd0;
            NN[254]=-25'd14;
            NN[255]=-25'd896;
            NN[256]=25'd1253;
            NN[257]=25'd14232;
            NN[258]=25'd18649;
            NN[259]=25'd12280;
            NN[260]=25'd3350;
            NN[261]=-25'd33;
            NN[262]=-25'd7259;
            NN[263]=-25'd12839;
            NN[264]=-25'd12720;
            NN[265]=-25'd15914;
            NN[266]=-25'd11224;
            NN[267]=25'd2144;
            NN[268]=25'd8058;
            NN[269]=25'd13982;
            NN[270]=25'd2744;
            NN[271]=-25'd489;
            NN[272]=-25'd3356;
            NN[273]=-25'd4782;
            NN[274]=-25'd3384;
            NN[275]=-25'd2462;
            NN[276]=-25'd625;
            NN[277]=-25'd77;
            NN[278]=25'd307;
            NN[279]=25'd0;
            NN[280]=25'd0;
            NN[281]=25'd0;
            NN[282]=25'd0;
            NN[283]=-25'd663;
            NN[284]=-25'd1096;
            NN[285]=25'd3244;
            NN[286]=25'd3623;
            NN[287]=-25'd2730;
            NN[288]=-25'd9085;
            NN[289]=-25'd11872;
            NN[290]=-25'd16705;
            NN[291]=-25'd20195;
            NN[292]=-25'd21901;
            NN[293]=-25'd24688;
            NN[294]=-25'd20803;
            NN[295]=-25'd15446;
            NN[296]=-25'd13198;
            NN[297]=-25'd4137;
            NN[298]=-25'd1745;
            NN[299]=-25'd525;
            NN[300]=-25'd1279;
            NN[301]=-25'd1005;
            NN[302]=-25'd1208;
            NN[303]=-25'd607;
            NN[304]=-25'd148;
            NN[305]=25'd192;
            NN[306]=25'd36;
            NN[307]=25'd0;
            NN[308]=25'd0;
            NN[309]=25'd0;
            NN[310]=25'd0;
            NN[311]=-25'd50;
            NN[312]=-25'd947;
            NN[313]=-25'd1756;
            NN[314]=-25'd2848;
            NN[315]=-25'd5349;
            NN[316]=-25'd6368;
            NN[317]=-25'd9488;
            NN[318]=-25'd14230;
            NN[319]=-25'd13823;
            NN[320]=-25'd12673;
            NN[321]=-25'd15750;
            NN[322]=-25'd15282;
            NN[323]=-25'd14537;
            NN[324]=-25'd10708;
            NN[325]=-25'd5454;
            NN[326]=-25'd1965;
            NN[327]=-25'd1348;
            NN[328]=-25'd634;
            NN[329]=-25'd229;
            NN[330]=-25'd159;
            NN[331]=-25'd26;
            NN[332]=25'd0;
            NN[333]=25'd0;
            NN[334]=25'd0;
            NN[335]=25'd0;
            NN[336]=25'd0;
            NN[337]=25'd0;
            NN[338]=25'd0;
            NN[339]=25'd0;
            NN[340]=-25'd59;
            NN[341]=-25'd136;
            NN[342]=-25'd229;
            NN[343]=-25'd427;
            NN[344]=-25'd790;
            NN[345]=-25'd1040;
            NN[346]=-25'd2092;
            NN[347]=-25'd1977;
            NN[348]=-25'd2578;
            NN[349]=-25'd4304;
            NN[350]=-25'd4057;
            NN[351]=-25'd3064;
            NN[352]=-25'd1813;
            NN[353]=-25'd710;
            NN[354]=-25'd425;
            NN[355]=-25'd204;
            NN[356]=-25'd101;
            NN[357]=-25'd60;
            NN[358]=-25'd15;
            NN[359]=-25'd1;
            NN[360]=25'd0;
            NN[361]=25'd0;
            NN[362]=25'd0;
            NN[363]=25'd0;
            NN[364]=25'd0;
            NN[365]=25'd0;
            NN[366]=25'd0;
            NN[367]=25'd0;
            NN[368]=25'd0;
            NN[369]=25'd0;
            NN[370]=25'd0;
            NN[371]=-25'd4;
            NN[372]=-25'd8;
            NN[373]=-25'd9;
            NN[374]=-25'd107;
            NN[375]=-25'd62;
            NN[376]=-25'd148;
            NN[377]=-25'd156;
            NN[378]=-25'd100;
            NN[379]=-25'd40;
            NN[380]=-25'd44;
            NN[381]=-25'd51;
            NN[382]=-25'd60;
            NN[383]=-25'd3;
            NN[384]=-25'd3;
            NN[385]=-25'd2;
            NN[386]=-25'd3;
            NN[387]=25'd0;
            NN[388]=25'd0;
            NN[389]=25'd0;
            NN[390]=25'd0;
            NN[391]=25'd0;
        end
        4:begin
            NN[0]=25'd0;
            NN[1]=25'd0;
            NN[2]=25'd0;
            NN[3]=25'd0;
            NN[4]=25'd0;
            NN[5]=25'd0;
            NN[6]=25'd0;
            NN[7]=25'd0;
            NN[8]=25'd0;
            NN[9]=25'd0;
            NN[10]=25'd0;
            NN[11]=25'd0;
            NN[12]=-25'd24;
            NN[13]=-25'd50;
            NN[14]=25'd2;
            NN[15]=25'd0;
            NN[16]=25'd0;
            NN[17]=25'd0;
            NN[18]=25'd0;
            NN[19]=25'd0;
            NN[20]=25'd0;
            NN[21]=25'd0;
            NN[22]=25'd0;
            NN[23]=25'd0;
            NN[24]=25'd0;
            NN[25]=25'd0;
            NN[26]=25'd0;
            NN[27]=25'd0;
            NN[28]=25'd0;
            NN[29]=25'd0;
            NN[30]=25'd0;
            NN[31]=25'd0;
            NN[32]=25'd0;
            NN[33]=-25'd1;
            NN[34]=-25'd14;
            NN[35]=-25'd33;
            NN[36]=-25'd110;
            NN[37]=-25'd240;
            NN[38]=-25'd403;
            NN[39]=-25'd472;
            NN[40]=-25'd656;
            NN[41]=-25'd397;
            NN[42]=25'd67;
            NN[43]=25'd337;
            NN[44]=25'd1319;
            NN[45]=25'd109;
            NN[46]=-25'd431;
            NN[47]=-25'd411;
            NN[48]=-25'd259;
            NN[49]=-25'd171;
            NN[50]=-25'd14;
            NN[51]=-25'd2;
            NN[52]=25'd0;
            NN[53]=25'd0;
            NN[54]=25'd0;
            NN[55]=25'd0;
            NN[56]=25'd0;
            NN[57]=25'd0;
            NN[58]=25'd0;
            NN[59]=25'd0;
            NN[60]=-25'd16;
            NN[61]=-25'd5;
            NN[62]=-25'd59;
            NN[63]=-25'd262;
            NN[64]=-25'd48;
            NN[65]=25'd1245;
            NN[66]=25'd395;
            NN[67]=25'd1904;
            NN[68]=25'd1106;
            NN[69]=25'd1032;
            NN[70]=25'd3039;
            NN[71]=25'd4500;
            NN[72]=25'd3705;
            NN[73]=25'd1339;
            NN[74]=-25'd923;
            NN[75]=-25'd2760;
            NN[76]=-25'd1778;
            NN[77]=-25'd1891;
            NN[78]=-25'd1798;
            NN[79]=-25'd676;
            NN[80]=25'd466;
            NN[81]=25'd415;
            NN[82]=25'd0;
            NN[83]=25'd0;
            NN[84]=25'd0;
            NN[85]=25'd0;
            NN[86]=25'd0;
            NN[87]=-25'd3;
            NN[88]=-25'd75;
            NN[89]=-25'd43;
            NN[90]=25'd80;
            NN[91]=25'd1248;
            NN[92]=25'd4147;
            NN[93]=25'd10314;
            NN[94]=25'd11544;
            NN[95]=25'd14194;
            NN[96]=25'd17069;
            NN[97]=25'd18256;
            NN[98]=25'd11246;
            NN[99]=25'd7518;
            NN[100]=25'd8385;
            NN[101]=25'd4156;
            NN[102]=-25'd4796;
            NN[103]=-25'd7814;
            NN[104]=-25'd9334;
            NN[105]=-25'd8247;
            NN[106]=-25'd6562;
            NN[107]=-25'd4185;
            NN[108]=-25'd1131;
            NN[109]=25'd207;
            NN[110]=-25'd17;
            NN[111]=25'd0;
            NN[112]=25'd0;
            NN[113]=25'd0;
            NN[114]=-25'd23;
            NN[115]=-25'd110;
            NN[116]=-25'd951;
            NN[117]=25'd168;
            NN[118]=25'd4065;
            NN[119]=25'd6501;
            NN[120]=25'd11591;
            NN[121]=25'd18908;
            NN[122]=25'd21564;
            NN[123]=25'd25342;
            NN[124]=25'd26542;
            NN[125]=25'd20497;
            NN[126]=25'd14869;
            NN[127]=25'd10247;
            NN[128]=25'd10777;
            NN[129]=25'd8608;
            NN[130]=25'd3945;
            NN[131]=-25'd4516;
            NN[132]=-25'd9100;
            NN[133]=-25'd13905;
            NN[134]=-25'd14463;
            NN[135]=-25'd9677;
            NN[136]=-25'd4850;
            NN[137]=-25'd677;
            NN[138]=-25'd84;
            NN[139]=-25'd59;
            NN[140]=25'd0;
            NN[141]=25'd0;
            NN[142]=25'd6;
            NN[143]=25'd87;
            NN[144]=-25'd260;
            NN[145]=25'd1103;
            NN[146]=25'd5586;
            NN[147]=25'd13405;
            NN[148]=25'd21301;
            NN[149]=25'd21601;
            NN[150]=25'd24084;
            NN[151]=25'd25167;
            NN[152]=25'd21750;
            NN[153]=25'd21393;
            NN[154]=25'd17643;
            NN[155]=25'd18299;
            NN[156]=25'd22328;
            NN[157]=25'd20452;
            NN[158]=25'd11448;
            NN[159]=25'd1025;
            NN[160]=-25'd3842;
            NN[161]=-25'd5503;
            NN[162]=-25'd10569;
            NN[163]=-25'd12631;
            NN[164]=-25'd8265;
            NN[165]=-25'd2182;
            NN[166]=-25'd340;
            NN[167]=-25'd86;
            NN[168]=25'd0;
            NN[169]=25'd0;
            NN[170]=-25'd109;
            NN[171]=25'd526;
            NN[172]=25'd1180;
            NN[173]=25'd4653;
            NN[174]=25'd12566;
            NN[175]=25'd18047;
            NN[176]=25'd17570;
            NN[177]=25'd18734;
            NN[178]=25'd14596;
            NN[179]=25'd6424;
            NN[180]=25'd7037;
            NN[181]=25'd8409;
            NN[182]=25'd9263;
            NN[183]=25'd8063;
            NN[184]=25'd8710;
            NN[185]=25'd5634;
            NN[186]=25'd2169;
            NN[187]=-25'd3693;
            NN[188]=-25'd7752;
            NN[189]=-25'd7286;
            NN[190]=-25'd10798;
            NN[191]=-25'd16251;
            NN[192]=-25'd9680;
            NN[193]=-25'd3177;
            NN[194]=-25'd353;
            NN[195]=-25'd19;
            NN[196]=25'd0;
            NN[197]=-25'd14;
            NN[198]=25'd279;
            NN[199]=25'd867;
            NN[200]=25'd5415;
            NN[201]=25'd8507;
            NN[202]=25'd16619;
            NN[203]=25'd12951;
            NN[204]=25'd13708;
            NN[205]=25'd7690;
            NN[206]=25'd2489;
            NN[207]=25'd5712;
            NN[208]=25'd1218;
            NN[209]=25'd5712;
            NN[210]=25'd3824;
            NN[211]=-25'd1862;
            NN[212]=-25'd4914;
            NN[213]=-25'd13032;
            NN[214]=-25'd8891;
            NN[215]=-25'd5457;
            NN[216]=-25'd6493;
            NN[217]=-25'd3116;
            NN[218]=-25'd2721;
            NN[219]=-25'd18450;
            NN[220]=-25'd13172;
            NN[221]=-25'd3881;
            NN[222]=-25'd465;
            NN[223]=-25'd29;
            NN[224]=-25'd1;
            NN[225]=25'd119;
            NN[226]=25'd197;
            NN[227]=25'd894;
            NN[228]=25'd6483;
            NN[229]=25'd9179;
            NN[230]=25'd10918;
            NN[231]=25'd9581;
            NN[232]=25'd8732;
            NN[233]=25'd8378;
            NN[234]=25'd17377;
            NN[235]=25'd13761;
            NN[236]=25'd6737;
            NN[237]=25'd3622;
            NN[238]=25'd7067;
            NN[239]=25'd3854;
            NN[240]=-25'd1918;
            NN[241]=-25'd3532;
            NN[242]=-25'd8207;
            NN[243]=25'd2177;
            NN[244]=-25'd2227;
            NN[245]=-25'd3246;
            NN[246]=-25'd4985;
            NN[247]=-25'd12541;
            NN[248]=-25'd14995;
            NN[249]=-25'd5584;
            NN[250]=-25'd582;
            NN[251]=-25'd28;
            NN[252]=25'd0;
            NN[253]=-25'd10;
            NN[254]=25'd45;
            NN[255]=25'd1546;
            NN[256]=25'd6377;
            NN[257]=25'd13097;
            NN[258]=25'd6172;
            NN[259]=25'd2147;
            NN[260]=-25'd1621;
            NN[261]=25'd7463;
            NN[262]=25'd14814;
            NN[263]=25'd9211;
            NN[264]=25'd5013;
            NN[265]=25'd6000;
            NN[266]=25'd10097;
            NN[267]=25'd11847;
            NN[268]=25'd12021;
            NN[269]=25'd5880;
            NN[270]=25'd6851;
            NN[271]=25'd1601;
            NN[272]=-25'd2590;
            NN[273]=-25'd5948;
            NN[274]=-25'd3110;
            NN[275]=-25'd11862;
            NN[276]=-25'd13696;
            NN[277]=-25'd4424;
            NN[278]=-25'd629;
            NN[279]=-25'd43;
            NN[280]=25'd0;
            NN[281]=-25'd5;
            NN[282]=25'd114;
            NN[283]=25'd2286;
            NN[284]=25'd558;
            NN[285]=25'd4814;
            NN[286]=25'd3214;
            NN[287]=-25'd10904;
            NN[288]=-25'd13166;
            NN[289]=-25'd12306;
            NN[290]=-25'd10181;
            NN[291]=-25'd13475;
            NN[292]=-25'd20162;
            NN[293]=-25'd23537;
            NN[294]=-25'd11999;
            NN[295]=-25'd5779;
            NN[296]=25'd1833;
            NN[297]=25'd4725;
            NN[298]=25'd7704;
            NN[299]=25'd392;
            NN[300]=-25'd2796;
            NN[301]=-25'd5666;
            NN[302]=-25'd4721;
            NN[303]=-25'd9564;
            NN[304]=-25'd8674;
            NN[305]=-25'd2473;
            NN[306]=-25'd234;
            NN[307]=-25'd21;
            NN[308]=25'd0;
            NN[309]=-25'd15;
            NN[310]=-25'd114;
            NN[311]=-25'd846;
            NN[312]=-25'd4695;
            NN[313]=-25'd10711;
            NN[314]=-25'd21011;
            NN[315]=-25'd32310;
            NN[316]=-25'd33868;
            NN[317]=-25'd37440;
            NN[318]=-25'd45684;
            NN[319]=-25'd47748;
            NN[320]=-25'd55434;
            NN[321]=-25'd54193;
            NN[322]=-25'd39331;
            NN[323]=-25'd27649;
            NN[324]=-25'd14112;
            NN[325]=-25'd15435;
            NN[326]=-25'd4758;
            NN[327]=25'd4450;
            NN[328]=-25'd2822;
            NN[329]=-25'd4409;
            NN[330]=-25'd8141;
            NN[331]=-25'd9905;
            NN[332]=-25'd4886;
            NN[333]=25'd440;
            NN[334]=25'd33;
            NN[335]=-25'd7;
            NN[336]=25'd0;
            NN[337]=-25'd3;
            NN[338]=-25'd21;
            NN[339]=-25'd2701;
            NN[340]=-25'd9415;
            NN[341]=-25'd26945;
            NN[342]=-25'd47896;
            NN[343]=-25'd54312;
            NN[344]=-25'd44878;
            NN[345]=-25'd46633;
            NN[346]=-25'd49875;
            NN[347]=-25'd49076;
            NN[348]=-25'd50517;
            NN[349]=-25'd43025;
            NN[350]=-25'd38279;
            NN[351]=-25'd32742;
            NN[352]=-25'd24834;
            NN[353]=-25'd22241;
            NN[354]=-25'd9780;
            NN[355]=25'd3844;
            NN[356]=-25'd1467;
            NN[357]=-25'd5537;
            NN[358]=-25'd11046;
            NN[359]=-25'd16736;
            NN[360]=-25'd1554;
            NN[361]=25'd5194;
            NN[362]=25'd2802;
            NN[363]=25'd318;
            NN[364]=25'd0;
            NN[365]=-25'd1;
            NN[366]=-25'd7;
            NN[367]=-25'd3002;
            NN[368]=-25'd13383;
            NN[369]=-25'd35151;
            NN[370]=-25'd52810;
            NN[371]=-25'd48940;
            NN[372]=-25'd36549;
            NN[373]=-25'd28773;
            NN[374]=-25'd20124;
            NN[375]=-25'd12243;
            NN[376]=-25'd12281;
            NN[377]=-25'd5459;
            NN[378]=-25'd9030;
            NN[379]=-25'd22423;
            NN[380]=-25'd24496;
            NN[381]=-25'd16833;
            NN[382]=-25'd13011;
            NN[383]=-25'd6636;
            NN[384]=-25'd6166;
            NN[385]=-25'd6000;
            NN[386]=-25'd11909;
            NN[387]=-25'd11951;
            NN[388]=25'd3294;
            NN[389]=25'd11442;
            NN[390]=25'd7188;
            NN[391]=25'd2041;
        end
        5:begin
            NN[0]=25'd0;
            NN[1]=-25'd160;
            NN[2]=-25'd110;
            NN[3]=-25'd2315;
            NN[4]=-25'd9335;
            NN[5]=-25'd27048;
            NN[6]=-25'd28615;
            NN[7]=-25'd18579;
            NN[8]=-25'd10372;
            NN[9]=-25'd2000;
            NN[10]=25'd4143;
            NN[11]=25'd9298;
            NN[12]=25'd8315;
            NN[13]=25'd19205;
            NN[14]=25'd5854;
            NN[15]=-25'd9264;
            NN[16]=-25'd8605;
            NN[17]=-25'd14713;
            NN[18]=-25'd8641;
            NN[19]=-25'd8201;
            NN[20]=-25'd3636;
            NN[21]=-25'd8423;
            NN[22]=-25'd11397;
            NN[23]=-25'd6075;
            NN[24]=25'd7215;
            NN[25]=25'd14541;
            NN[26]=25'd7840;
            NN[27]=25'd335;
            NN[28]=25'd0;
            NN[29]=-25'd344;
            NN[30]=-25'd94;
            NN[31]=25'd1254;
            NN[32]=25'd1488;
            NN[33]=-25'd1866;
            NN[34]=25'd985;
            NN[35]=25'd1619;
            NN[36]=25'd2071;
            NN[37]=25'd5616;
            NN[38]=25'd3870;
            NN[39]=25'd640;
            NN[40]=25'd9836;
            NN[41]=25'd18630;
            NN[42]=25'd8199;
            NN[43]=25'd656;
            NN[44]=-25'd647;
            NN[45]=-25'd7781;
            NN[46]=-25'd13336;
            NN[47]=-25'd6315;
            NN[48]=-25'd12507;
            NN[49]=-25'd10535;
            NN[50]=-25'd12382;
            NN[51]=-25'd2271;
            NN[52]=25'd17879;
            NN[53]=25'd21688;
            NN[54]=25'd9626;
            NN[55]=25'd1289;
            NN[56]=25'd0;
            NN[57]=-25'd178;
            NN[58]=25'd105;
            NN[59]=25'd5651;
            NN[60]=25'd12095;
            NN[61]=25'd12323;
            NN[62]=25'd16826;
            NN[63]=25'd8239;
            NN[64]=25'd1945;
            NN[65]=25'd8803;
            NN[66]=25'd8028;
            NN[67]=25'd14633;
            NN[68]=25'd21837;
            NN[69]=25'd25454;
            NN[70]=25'd11050;
            NN[71]=25'd1883;
            NN[72]=25'd11846;
            NN[73]=25'd7965;
            NN[74]=-25'd176;
            NN[75]=-25'd1668;
            NN[76]=-25'd3060;
            NN[77]=25'd8898;
            NN[78]=25'd9240;
            NN[79]=25'd13500;
            NN[80]=25'd27260;
            NN[81]=25'd32430;
            NN[82]=25'd12775;
            NN[83]=25'd1363;
            NN[84]=25'd0;
            NN[85]=-25'd72;
            NN[86]=25'd727;
            NN[87]=25'd8154;
            NN[88]=25'd21678;
            NN[89]=25'd23524;
            NN[90]=25'd19554;
            NN[91]=25'd13325;
            NN[92]=25'd11457;
            NN[93]=25'd12419;
            NN[94]=25'd16470;
            NN[95]=25'd22001;
            NN[96]=25'd29854;
            NN[97]=25'd23535;
            NN[98]=25'd8673;
            NN[99]=25'd9400;
            NN[100]=25'd9573;
            NN[101]=25'd4135;
            NN[102]=25'd3012;
            NN[103]=25'd1203;
            NN[104]=25'd4726;
            NN[105]=25'd12499;
            NN[106]=25'd17319;
            NN[107]=25'd19608;
            NN[108]=25'd34885;
            NN[109]=25'd34662;
            NN[110]=25'd8069;
            NN[111]=25'd560;
            NN[112]=-25'd3;
            NN[113]=-25'd8;
            NN[114]=-25'd452;
            NN[115]=25'd6884;
            NN[116]=25'd23732;
            NN[117]=25'd29451;
            NN[118]=25'd19683;
            NN[119]=25'd23267;
            NN[120]=25'd12605;
            NN[121]=25'd13048;
            NN[122]=25'd18154;
            NN[123]=25'd18433;
            NN[124]=25'd25530;
            NN[125]=25'd24260;
            NN[126]=25'd14304;
            NN[127]=25'd4674;
            NN[128]=25'd9988;
            NN[129]=25'd11817;
            NN[130]=25'd8295;
            NN[131]=25'd7227;
            NN[132]=25'd6520;
            NN[133]=25'd13360;
            NN[134]=25'd18266;
            NN[135]=25'd32159;
            NN[136]=25'd40932;
            NN[137]=25'd25055;
            NN[138]=25'd2917;
            NN[139]=25'd896;
            NN[140]=25'd0;
            NN[141]=-25'd65;
            NN[142]=-25'd348;
            NN[143]=25'd2596;
            NN[144]=25'd18022;
            NN[145]=25'd20284;
            NN[146]=25'd19703;
            NN[147]=25'd25325;
            NN[148]=25'd20934;
            NN[149]=25'd20369;
            NN[150]=25'd22657;
            NN[151]=25'd22315;
            NN[152]=25'd22182;
            NN[153]=25'd25166;
            NN[154]=25'd12603;
            NN[155]=25'd8111;
            NN[156]=25'd7936;
            NN[157]=25'd10456;
            NN[158]=25'd7148;
            NN[159]=25'd4590;
            NN[160]=25'd9643;
            NN[161]=25'd17708;
            NN[162]=25'd26712;
            NN[163]=25'd30652;
            NN[164]=25'd28298;
            NN[165]=25'd16621;
            NN[166]=25'd3951;
            NN[167]=25'd455;
            NN[168]=25'd0;
            NN[169]=-25'd144;
            NN[170]=-25'd31;
            NN[171]=25'd3769;
            NN[172]=25'd15969;
            NN[173]=25'd17943;
            NN[174]=25'd18907;
            NN[175]=25'd28089;
            NN[176]=25'd23576;
            NN[177]=25'd20062;
            NN[178]=25'd15170;
            NN[179]=25'd17583;
            NN[180]=25'd11394;
            NN[181]=25'd5236;
            NN[182]=25'd1398;
            NN[183]=25'd1438;
            NN[184]=25'd3669;
            NN[185]=25'd3535;
            NN[186]=25'd10739;
            NN[187]=25'd13318;
            NN[188]=25'd12100;
            NN[189]=25'd20499;
            NN[190]=25'd27792;
            NN[191]=25'd28159;
            NN[192]=25'd22905;
            NN[193]=25'd7911;
            NN[194]=25'd1562;
            NN[195]=-25'd4;
            NN[196]=25'd0;
            NN[197]=25'd2;
            NN[198]=25'd13;
            NN[199]=25'd2738;
            NN[200]=25'd8841;
            NN[201]=25'd10857;
            NN[202]=25'd13957;
            NN[203]=25'd15177;
            NN[204]=25'd14753;
            NN[205]=25'd18981;
            NN[206]=25'd12166;
            NN[207]=25'd9151;
            NN[208]=25'd2480;
            NN[209]=25'd4024;
            NN[210]=-25'd107;
            NN[211]=-25'd2816;
            NN[212]=25'd4462;
            NN[213]=25'd10045;
            NN[214]=25'd15579;
            NN[215]=25'd20434;
            NN[216]=25'd12037;
            NN[217]=25'd19294;
            NN[218]=25'd26413;
            NN[219]=25'd25990;
            NN[220]=25'd15925;
            NN[221]=25'd4902;
            NN[222]=25'd750;
            NN[223]=25'd0;
            NN[224]=25'd0;
            NN[225]=25'd0;
            NN[226]=25'd78;
            NN[227]=25'd1383;
            NN[228]=25'd5005;
            NN[229]=25'd5347;
            NN[230]=25'd10442;
            NN[231]=25'd12727;
            NN[232]=25'd18362;
            NN[233]=25'd19184;
            NN[234]=25'd14179;
            NN[235]=25'd10235;
            NN[236]=25'd5647;
            NN[237]=-25'd1957;
            NN[238]=-25'd8281;
            NN[239]=-25'd10800;
            NN[240]=-25'd3565;
            NN[241]=25'd1669;
            NN[242]=25'd13537;
            NN[243]=25'd19693;
            NN[244]=25'd18777;
            NN[245]=25'd20324;
            NN[246]=25'd19844;
            NN[247]=25'd13179;
            NN[248]=25'd7303;
            NN[249]=25'd1722;
            NN[250]=-25'd365;
            NN[251]=25'd0;
            NN[252]=25'd0;
            NN[253]=25'd0;
            NN[254]=-25'd104;
            NN[255]=-25'd795;
            NN[256]=-25'd1252;
            NN[257]=-25'd3236;
            NN[258]=-25'd3912;
            NN[259]=-25'd3666;
            NN[260]=25'd494;
            NN[261]=25'd2175;
            NN[262]=25'd777;
            NN[263]=25'd3630;
            NN[264]=-25'd1840;
            NN[265]=-25'd12981;
            NN[266]=-25'd15696;
            NN[267]=-25'd14199;
            NN[268]=-25'd7976;
            NN[269]=-25'd2735;
            NN[270]=25'd9321;
            NN[271]=25'd14892;
            NN[272]=25'd10919;
            NN[273]=25'd13631;
            NN[274]=25'd10760;
            NN[275]=25'd5535;
            NN[276]=25'd3680;
            NN[277]=25'd1314;
            NN[278]=-25'd263;
            NN[279]=25'd0;
            NN[280]=25'd0;
            NN[281]=25'd0;
            NN[282]=-25'd79;
            NN[283]=-25'd1654;
            NN[284]=-25'd3804;
            NN[285]=-25'd8073;
            NN[286]=-25'd13007;
            NN[287]=-25'd17865;
            NN[288]=-25'd17777;
            NN[289]=-25'd17282;
            NN[290]=-25'd20454;
            NN[291]=-25'd15396;
            NN[292]=-25'd9319;
            NN[293]=-25'd7811;
            NN[294]=-25'd3077;
            NN[295]=-25'd6311;
            NN[296]=-25'd4480;
            NN[297]=-25'd947;
            NN[298]=25'd284;
            NN[299]=-25'd5684;
            NN[300]=-25'd3378;
            NN[301]=25'd1493;
            NN[302]=25'd1540;
            NN[303]=25'd1541;
            NN[304]=25'd4072;
            NN[305]=25'd2275;
            NN[306]=25'd321;
            NN[307]=25'd0;
            NN[308]=25'd0;
            NN[309]=25'd0;
            NN[310]=-25'd1;
            NN[311]=-25'd381;
            NN[312]=-25'd1570;
            NN[313]=-25'd2788;
            NN[314]=-25'd4052;
            NN[315]=-25'd8333;
            NN[316]=-25'd13926;
            NN[317]=-25'd14321;
            NN[318]=-25'd11850;
            NN[319]=-25'd10881;
            NN[320]=-25'd9418;
            NN[321]=-25'd8410;
            NN[322]=-25'd5985;
            NN[323]=-25'd4280;
            NN[324]=-25'd3889;
            NN[325]=-25'd4354;
            NN[326]=-25'd6713;
            NN[327]=-25'd8148;
            NN[328]=-25'd4821;
            NN[329]=-25'd3548;
            NN[330]=-25'd2462;
            NN[331]=-25'd1315;
            NN[332]=-25'd142;
            NN[333]=25'd284;
            NN[334]=25'd341;
            NN[335]=25'd0;
            NN[336]=25'd0;
            NN[337]=25'd0;
            NN[338]=25'd0;
            NN[339]=25'd0;
            NN[340]=-25'd59;
            NN[341]=-25'd170;
            NN[342]=-25'd379;
            NN[343]=-25'd891;
            NN[344]=-25'd984;
            NN[345]=-25'd846;
            NN[346]=-25'd907;
            NN[347]=-25'd1515;
            NN[348]=-25'd1290;
            NN[349]=-25'd1724;
            NN[350]=-25'd1432;
            NN[351]=-25'd1486;
            NN[352]=-25'd1726;
            NN[353]=-25'd1763;
            NN[354]=-25'd1587;
            NN[355]=-25'd1049;
            NN[356]=-25'd601;
            NN[357]=-25'd553;
            NN[358]=-25'd180;
            NN[359]=-25'd3;
            NN[360]=25'd0;
            NN[361]=25'd0;
            NN[362]=25'd0;
            NN[363]=25'd0;
            NN[364]=25'd0;
            NN[365]=25'd0;
            NN[366]=25'd0;
            NN[367]=25'd0;
            NN[368]=25'd0;
            NN[369]=25'd0;
            NN[370]=-25'd1;
            NN[371]=-25'd20;
            NN[372]=-25'd27;
            NN[373]=-25'd28;
            NN[374]=-25'd48;
            NN[375]=-25'd44;
            NN[376]=-25'd45;
            NN[377]=-25'd57;
            NN[378]=-25'd97;
            NN[379]=-25'd94;
            NN[380]=-25'd112;
            NN[381]=-25'd118;
            NN[382]=-25'd22;
            NN[383]=-25'd7;
            NN[384]=-25'd47;
            NN[385]=-25'd39;
            NN[386]=-25'd166;
            NN[387]=-25'd3;
            NN[388]=25'd0;
            NN[389]=25'd0;
            NN[390]=25'd0;
            NN[391]=25'd0;
        end
        6:begin
            NN[0]=25'd0;
            NN[1]=25'd0;
            NN[2]=25'd0;
            NN[3]=25'd0;
            NN[4]=25'd0;
            NN[5]=25'd0;
            NN[6]=25'd0;
            NN[7]=25'd0;
            NN[8]=25'd0;
            NN[9]=25'd0;
            NN[10]=25'd0;
            NN[11]=25'd0;
            NN[12]=-25'd1;
            NN[13]=-25'd2;
            NN[14]=25'd0;
            NN[15]=25'd0;
            NN[16]=25'd0;
            NN[17]=25'd0;
            NN[18]=25'd0;
            NN[19]=25'd0;
            NN[20]=25'd0;
            NN[21]=25'd0;
            NN[22]=25'd0;
            NN[23]=25'd0;
            NN[24]=25'd0;
            NN[25]=25'd0;
            NN[26]=25'd0;
            NN[27]=25'd0;
            NN[28]=25'd0;
            NN[29]=25'd0;
            NN[30]=25'd0;
            NN[31]=25'd0;
            NN[32]=25'd0;
            NN[33]=25'd0;
            NN[34]=25'd0;
            NN[35]=25'd0;
            NN[36]=-25'd8;
            NN[37]=-25'd42;
            NN[38]=-25'd120;
            NN[39]=-25'd53;
            NN[40]=-25'd95;
            NN[41]=-25'd123;
            NN[42]=-25'd83;
            NN[43]=-25'd75;
            NN[44]=-25'd77;
            NN[45]=-25'd25;
            NN[46]=-25'd6;
            NN[47]=-25'd6;
            NN[48]=-25'd8;
            NN[49]=-25'd2;
            NN[50]=25'd0;
            NN[51]=25'd0;
            NN[52]=25'd0;
            NN[53]=25'd0;
            NN[54]=25'd0;
            NN[55]=25'd0;
            NN[56]=25'd0;
            NN[57]=25'd0;
            NN[58]=25'd0;
            NN[59]=25'd0;
            NN[60]=25'd0;
            NN[61]=-25'd2;
            NN[62]=-25'd17;
            NN[63]=-25'd81;
            NN[64]=-25'd262;
            NN[65]=-25'd688;
            NN[66]=-25'd637;
            NN[67]=25'd69;
            NN[68]=25'd208;
            NN[69]=-25'd142;
            NN[70]=25'd76;
            NN[71]=-25'd548;
            NN[72]=-25'd601;
            NN[73]=-25'd357;
            NN[74]=-25'd290;
            NN[75]=-25'd332;
            NN[76]=-25'd395;
            NN[77]=-25'd438;
            NN[78]=-25'd341;
            NN[79]=-25'd78;
            NN[80]=-25'd11;
            NN[81]=25'd0;
            NN[82]=25'd0;
            NN[83]=25'd0;
            NN[84]=25'd0;
            NN[85]=25'd0;
            NN[86]=25'd0;
            NN[87]=-25'd1;
            NN[88]=-25'd42;
            NN[89]=25'd1319;
            NN[90]=25'd1150;
            NN[91]=25'd2062;
            NN[92]=25'd2662;
            NN[93]=25'd2107;
            NN[94]=25'd5252;
            NN[95]=25'd11233;
            NN[96]=25'd15525;
            NN[97]=25'd14543;
            NN[98]=25'd19905;
            NN[99]=25'd19943;
            NN[100]=25'd16587;
            NN[101]=25'd14187;
            NN[102]=25'd11995;
            NN[103]=25'd8407;
            NN[104]=25'd5242;
            NN[105]=-25'd1416;
            NN[106]=-25'd2685;
            NN[107]=-25'd1266;
            NN[108]=-25'd452;
            NN[109]=-25'd37;
            NN[110]=25'd0;
            NN[111]=25'd0;
            NN[112]=25'd0;
            NN[113]=25'd1;
            NN[114]=25'd39;
            NN[115]=25'd384;
            NN[116]=25'd1790;
            NN[117]=25'd6328;
            NN[118]=25'd9052;
            NN[119]=25'd12606;
            NN[120]=25'd17645;
            NN[121]=25'd20602;
            NN[122]=25'd23624;
            NN[123]=25'd28133;
            NN[124]=25'd26899;
            NN[125]=25'd26667;
            NN[126]=25'd23604;
            NN[127]=25'd22007;
            NN[128]=25'd21211;
            NN[129]=25'd13484;
            NN[130]=25'd11820;
            NN[131]=25'd3696;
            NN[132]=-25'd5006;
            NN[133]=-25'd8958;
            NN[134]=-25'd7601;
            NN[135]=-25'd7747;
            NN[136]=-25'd1938;
            NN[137]=-25'd237;
            NN[138]=-25'd45;
            NN[139]=-25'd2;
            NN[140]=25'd0;
            NN[141]=25'd0;
            NN[142]=25'd147;
            NN[143]=25'd2054;
            NN[144]=25'd5929;
            NN[145]=25'd14073;
            NN[146]=25'd19240;
            NN[147]=25'd20092;
            NN[148]=25'd18954;
            NN[149]=25'd20561;
            NN[150]=25'd18747;
            NN[151]=25'd14744;
            NN[152]=25'd10468;
            NN[153]=25'd8493;
            NN[154]=25'd5803;
            NN[155]=25'd11366;
            NN[156]=25'd14429;
            NN[157]=25'd586;
            NN[158]=-25'd528;
            NN[159]=-25'd424;
            NN[160]=-25'd6182;
            NN[161]=-25'd12560;
            NN[162]=-25'd14236;
            NN[163]=-25'd13616;
            NN[164]=-25'd5310;
            NN[165]=-25'd1130;
            NN[166]=-25'd142;
            NN[167]=-25'd6;
            NN[168]=25'd0;
            NN[169]=25'd6;
            NN[170]=25'd318;
            NN[171]=25'd4108;
            NN[172]=25'd10138;
            NN[173]=25'd16848;
            NN[174]=25'd19685;
            NN[175]=25'd14965;
            NN[176]=25'd16344;
            NN[177]=25'd20100;
            NN[178]=25'd17452;
            NN[179]=25'd11394;
            NN[180]=25'd10953;
            NN[181]=25'd17194;
            NN[182]=25'd12445;
            NN[183]=25'd13754;
            NN[184]=25'd17288;
            NN[185]=25'd11253;
            NN[186]=25'd12146;
            NN[187]=-25'd967;
            NN[188]=25'd2386;
            NN[189]=-25'd2280;
            NN[190]=-25'd12893;
            NN[191]=-25'd15591;
            NN[192]=-25'd7176;
            NN[193]=-25'd2227;
            NN[194]=-25'd324;
            NN[195]=-25'd9;
            NN[196]=25'd0;
            NN[197]=25'd200;
            NN[198]=25'd213;
            NN[199]=25'd4274;
            NN[200]=25'd15448;
            NN[201]=25'd21120;
            NN[202]=25'd17734;
            NN[203]=25'd10829;
            NN[204]=25'd7660;
            NN[205]=25'd6314;
            NN[206]=25'd4951;
            NN[207]=25'd4303;
            NN[208]=25'd9951;
            NN[209]=25'd12042;
            NN[210]=25'd17767;
            NN[211]=25'd19861;
            NN[212]=25'd10352;
            NN[213]=25'd10648;
            NN[214]=25'd5981;
            NN[215]=25'd8754;
            NN[216]=25'd6985;
            NN[217]=25'd788;
            NN[218]=-25'd9972;
            NN[219]=-25'd16602;
            NN[220]=-25'd11099;
            NN[221]=-25'd2984;
            NN[222]=-25'd272;
            NN[223]=-25'd14;
            NN[224]=25'd0;
            NN[225]=-25'd94;
            NN[226]=25'd101;
            NN[227]=25'd4284;
            NN[228]=25'd15644;
            NN[229]=25'd16536;
            NN[230]=25'd12786;
            NN[231]=25'd8782;
            NN[232]=25'd5419;
            NN[233]=25'd2851;
            NN[234]=25'd5264;
            NN[235]=-25'd1309;
            NN[236]=25'd1380;
            NN[237]=25'd8432;
            NN[238]=25'd20180;
            NN[239]=25'd24223;
            NN[240]=25'd15824;
            NN[241]=25'd13205;
            NN[242]=25'd12730;
            NN[243]=25'd13013;
            NN[244]=25'd14872;
            NN[245]=25'd12428;
            NN[246]=25'd1818;
            NN[247]=-25'd19577;
            NN[248]=-25'd14325;
            NN[249]=-25'd3593;
            NN[250]=-25'd311;
            NN[251]=-25'd4;
            NN[252]=-25'd4;
            NN[253]=-25'd91;
            NN[254]=25'd529;
            NN[255]=25'd4798;
            NN[256]=25'd15366;
            NN[257]=25'd10290;
            NN[258]=25'd8657;
            NN[259]=25'd2877;
            NN[260]=-25'd4450;
            NN[261]=-25'd8606;
            NN[262]=-25'd17945;
            NN[263]=-25'd32213;
            NN[264]=-25'd24959;
            NN[265]=-25'd7139;
            NN[266]=25'd17892;
            NN[267]=25'd27685;
            NN[268]=25'd22394;
            NN[269]=25'd14157;
            NN[270]=25'd9430;
            NN[271]=25'd15701;
            NN[272]=25'd23791;
            NN[273]=25'd17516;
            NN[274]=25'd4759;
            NN[275]=-25'd12668;
            NN[276]=-25'd11954;
            NN[277]=-25'd2623;
            NN[278]=-25'd462;
            NN[279]=-25'd13;
            NN[280]=-25'd5;
            NN[281]=-25'd85;
            NN[282]=25'd331;
            NN[283]=25'd5886;
            NN[284]=25'd7352;
            NN[285]=25'd1262;
            NN[286]=-25'd6406;
            NN[287]=-25'd16161;
            NN[288]=-25'd25837;
            NN[289]=-25'd35797;
            NN[290]=-25'd42017;
            NN[291]=-25'd45066;
            NN[292]=-25'd33774;
            NN[293]=25'd53;
            NN[294]=25'd21297;
            NN[295]=25'd20686;
            NN[296]=25'd21524;
            NN[297]=25'd15247;
            NN[298]=25'd14459;
            NN[299]=25'd19856;
            NN[300]=25'd22771;
            NN[301]=25'd10332;
            NN[302]=-25'd413;
            NN[303]=-25'd8022;
            NN[304]=-25'd7553;
            NN[305]=-25'd1446;
            NN[306]=-25'd249;
            NN[307]=-25'd4;
            NN[308]=-25'd4;
            NN[309]=-25'd106;
            NN[310]=25'd75;
            NN[311]=25'd5084;
            NN[312]=25'd2159;
            NN[313]=-25'd9093;
            NN[314]=-25'd20897;
            NN[315]=-25'd33744;
            NN[316]=-25'd37377;
            NN[317]=-25'd35563;
            NN[318]=-25'd29047;
            NN[319]=-25'd20648;
            NN[320]=-25'd6670;
            NN[321]=25'd13627;
            NN[322]=25'd18336;
            NN[323]=25'd19613;
            NN[324]=25'd11394;
            NN[325]=25'd16912;
            NN[326]=25'd15839;
            NN[327]=25'd17630;
            NN[328]=25'd13368;
            NN[329]=-25'd5409;
            NN[330]=-25'd8203;
            NN[331]=-25'd8402;
            NN[332]=-25'd5421;
            NN[333]=-25'd507;
            NN[334]=-25'd84;
            NN[335]=-25'd1;
            NN[336]=-25'd2;
            NN[337]=-25'd142;
            NN[338]=-25'd620;
            NN[339]=25'd456;
            NN[340]=-25'd3091;
            NN[341]=-25'd14049;
            NN[342]=-25'd24802;
            NN[343]=-25'd32415;
            NN[344]=-25'd31068;
            NN[345]=-25'd17767;
            NN[346]=-25'd4126;
            NN[347]=-25'd6674;
            NN[348]=25'd3200;
            NN[349]=25'd13331;
            NN[350]=25'd27380;
            NN[351]=25'd17234;
            NN[352]=25'd11842;
            NN[353]=25'd13637;
            NN[354]=25'd13417;
            NN[355]=25'd1223;
            NN[356]=-25'd8618;
            NN[357]=-25'd21535;
            NN[358]=-25'd15938;
            NN[359]=-25'd9341;
            NN[360]=-25'd4014;
            NN[361]=25'd14;
            NN[362]=-25'd18;
            NN[363]=-25'd2;
            NN[364]=25'd0;
            NN[365]=-25'd94;
            NN[366]=-25'd473;
            NN[367]=-25'd499;
            NN[368]=-25'd6016;
            NN[369]=-25'd14877;
            NN[370]=-25'd23353;
            NN[371]=-25'd28828;
            NN[372]=-25'd21706;
            NN[373]=-25'd11395;
            NN[374]=-25'd14695;
            NN[375]=-25'd13305;
            NN[376]=25'd6281;
            NN[377]=25'd20008;
            NN[378]=25'd17352;
            NN[379]=25'd660;
            NN[380]=25'd9922;
            NN[381]=25'd12017;
            NN[382]=25'd9745;
            NN[383]=-25'd6644;
            NN[384]=-25'd21917;
            NN[385]=-25'd20870;
            NN[386]=-25'd19072;
            NN[387]=-25'd9636;
            NN[388]=-25'd3658;
            NN[389]=-25'd348;
            NN[390]=-25'd63;
            NN[391]=-25'd86;
        end
        7:begin
            NN[0]=-25'd68;
            NN[1]=25'd232;
            NN[2]=-25'd8;
            NN[3]=25'd190;
            NN[4]=-25'd3016;
            NN[5]=-25'd13322;
            NN[6]=-25'd22770;
            NN[7]=-25'd24921;
            NN[8]=-25'd19080;
            NN[9]=-25'd16286;
            NN[10]=-25'd19458;
            NN[11]=-25'd16579;
            NN[12]=25'd6876;
            NN[13]=25'd10107;
            NN[14]=25'd10870;
            NN[15]=25'd3788;
            NN[16]=25'd4218;
            NN[17]=25'd7828;
            NN[18]=25'd4701;
            NN[19]=-25'd3931;
            NN[20]=-25'd10037;
            NN[21]=-25'd4000;
            NN[22]=-25'd11983;
            NN[23]=-25'd8301;
            NN[24]=-25'd2750;
            NN[25]=-25'd970;
            NN[26]=-25'd459;
            NN[27]=-25'd70;
            NN[28]=-25'd22;
            NN[29]=25'd592;
            NN[30]=25'd597;
            NN[31]=25'd1658;
            NN[32]=25'd1849;
            NN[33]=-25'd6025;
            NN[34]=-25'd13549;
            NN[35]=-25'd19585;
            NN[36]=-25'd23479;
            NN[37]=-25'd25717;
            NN[38]=-25'd20278;
            NN[39]=-25'd8369;
            NN[40]=25'd4157;
            NN[41]=25'd11999;
            NN[42]=25'd10883;
            NN[43]=-25'd332;
            NN[44]=-25'd5972;
            NN[45]=25'd1603;
            NN[46]=25'd3593;
            NN[47]=25'd9227;
            NN[48]=25'd14070;
            NN[49]=25'd12267;
            NN[50]=25'd6571;
            NN[51]=25'd1536;
            NN[52]=-25'd315;
            NN[53]=-25'd1810;
            NN[54]=-25'd617;
            NN[55]=-25'd46;
            NN[56]=25'd0;
            NN[57]=25'd406;
            NN[58]=25'd1871;
            NN[59]=25'd5723;
            NN[60]=25'd9773;
            NN[61]=25'd2516;
            NN[62]=-25'd8403;
            NN[63]=-25'd15061;
            NN[64]=-25'd24148;
            NN[65]=-25'd23539;
            NN[66]=-25'd23668;
            NN[67]=-25'd11959;
            NN[68]=-25'd117;
            NN[69]=25'd9106;
            NN[70]=-25'd4633;
            NN[71]=-25'd17768;
            NN[72]=-25'd16019;
            NN[73]=25'd529;
            NN[74]=25'd16250;
            NN[75]=25'd19744;
            NN[76]=25'd17076;
            NN[77]=25'd18926;
            NN[78]=25'd18066;
            NN[79]=25'd10440;
            NN[80]=25'd2988;
            NN[81]=-25'd2678;
            NN[82]=-25'd578;
            NN[83]=-25'd30;
            NN[84]=25'd0;
            NN[85]=25'd121;
            NN[86]=25'd2394;
            NN[87]=25'd11636;
            NN[88]=25'd15803;
            NN[89]=25'd6632;
            NN[90]=-25'd4486;
            NN[91]=-25'd10821;
            NN[92]=-25'd21970;
            NN[93]=-25'd36625;
            NN[94]=-25'd41310;
            NN[95]=-25'd34429;
            NN[96]=-25'd26696;
            NN[97]=-25'd21925;
            NN[98]=-25'd23803;
            NN[99]=-25'd18838;
            NN[100]=-25'd565;
            NN[101]=25'd12562;
            NN[102]=25'd12525;
            NN[103]=25'd20000;
            NN[104]=25'd14332;
            NN[105]=25'd21830;
            NN[106]=25'd24553;
            NN[107]=25'd13968;
            NN[108]=-25'd3208;
            NN[109]=-25'd4463;
            NN[110]=-25'd490;
            NN[111]=-25'd18;
            NN[112]=-25'd19;
            NN[113]=25'd16;
            NN[114]=25'd2636;
            NN[115]=25'd17957;
            NN[116]=25'd21461;
            NN[117]=25'd17215;
            NN[118]=25'd6807;
            NN[119]=-25'd6740;
            NN[120]=-25'd14643;
            NN[121]=-25'd28127;
            NN[122]=-25'd36024;
            NN[123]=-25'd36904;
            NN[124]=-25'd37004;
            NN[125]=-25'd30738;
            NN[126]=-25'd24808;
            NN[127]=-25'd938;
            NN[128]=25'd19756;
            NN[129]=25'd18405;
            NN[130]=25'd18022;
            NN[131]=25'd16943;
            NN[132]=25'd14447;
            NN[133]=25'd27406;
            NN[134]=25'd26873;
            NN[135]=25'd7972;
            NN[136]=-25'd7383;
            NN[137]=-25'd3725;
            NN[138]=-25'd538;
            NN[139]=-25'd19;
            NN[140]=25'd0;
            NN[141]=-25'd7;
            NN[142]=25'd2794;
            NN[143]=25'd22042;
            NN[144]=25'd25798;
            NN[145]=25'd24523;
            NN[146]=25'd13157;
            NN[147]=25'd5721;
            NN[148]=25'd1534;
            NN[149]=-25'd5885;
            NN[150]=-25'd15315;
            NN[151]=-25'd22175;
            NN[152]=-25'd24942;
            NN[153]=-25'd20006;
            NN[154]=-25'd12491;
            NN[155]=25'd2486;
            NN[156]=25'd16033;
            NN[157]=25'd21777;
            NN[158]=25'd24005;
            NN[159]=25'd17660;
            NN[160]=25'd16774;
            NN[161]=25'd24062;
            NN[162]=25'd12774;
            NN[163]=25'd2585;
            NN[164]=-25'd6157;
            NN[165]=-25'd2522;
            NN[166]=-25'd475;
            NN[167]=-25'd13;
            NN[168]=25'd0;
            NN[169]=-25'd21;
            NN[170]=25'd2637;
            NN[171]=25'd19801;
            NN[172]=25'd26731;
            NN[173]=25'd23143;
            NN[174]=25'd21196;
            NN[175]=25'd15909;
            NN[176]=25'd15141;
            NN[177]=25'd13661;
            NN[178]=-25'd570;
            NN[179]=-25'd12917;
            NN[180]=-25'd19767;
            NN[181]=-25'd10149;
            NN[182]=-25'd816;
            NN[183]=25'd2327;
            NN[184]=25'd11469;
            NN[185]=25'd17048;
            NN[186]=25'd22188;
            NN[187]=25'd17157;
            NN[188]=25'd22337;
            NN[189]=25'd11961;
            NN[190]=25'd131;
            NN[191]=-25'd3030;
            NN[192]=-25'd5439;
            NN[193]=-25'd1395;
            NN[194]=-25'd181;
            NN[195]=25'd0;
            NN[196]=25'd0;
            NN[197]=25'd21;
            NN[198]=25'd3155;
            NN[199]=25'd13439;
            NN[200]=25'd20294;
            NN[201]=25'd18440;
            NN[202]=25'd18760;
            NN[203]=25'd12595;
            NN[204]=25'd8590;
            NN[205]=25'd1126;
            NN[206]=-25'd1743;
            NN[207]=-25'd7741;
            NN[208]=-25'd7940;
            NN[209]=-25'd4001;
            NN[210]=-25'd1875;
            NN[211]=25'd3328;
            NN[212]=25'd9037;
            NN[213]=25'd8620;
            NN[214]=25'd16964;
            NN[215]=25'd18382;
            NN[216]=25'd9500;
            NN[217]=-25'd2942;
            NN[218]=-25'd6832;
            NN[219]=-25'd8325;
            NN[220]=-25'd5594;
            NN[221]=-25'd1385;
            NN[222]=-25'd228;
            NN[223]=25'd0;
            NN[224]=25'd0;
            NN[225]=25'd0;
            NN[226]=25'd3084;
            NN[227]=25'd9057;
            NN[228]=25'd14111;
            NN[229]=25'd16263;
            NN[230]=25'd17214;
            NN[231]=25'd9088;
            NN[232]=-25'd2455;
            NN[233]=25'd677;
            NN[234]=25'd2522;
            NN[235]=25'd2499;
            NN[236]=-25'd5176;
            NN[237]=-25'd4200;
            NN[238]=-25'd1704;
            NN[239]=25'd2696;
            NN[240]=25'd4024;
            NN[241]=25'd6272;
            NN[242]=25'd10520;
            NN[243]=25'd11238;
            NN[244]=25'd3204;
            NN[245]=-25'd6085;
            NN[246]=-25'd4029;
            NN[247]=-25'd4972;
            NN[248]=-25'd3113;
            NN[249]=-25'd777;
            NN[250]=-25'd11;
            NN[251]=25'd0;
            NN[252]=25'd0;
            NN[253]=25'd0;
            NN[254]=25'd1430;
            NN[255]=25'd6195;
            NN[256]=25'd12836;
            NN[257]=25'd19924;
            NN[258]=25'd21764;
            NN[259]=25'd17784;
            NN[260]=25'd5341;
            NN[261]=25'd6058;
            NN[262]=25'd6126;
            NN[263]=25'd7671;
            NN[264]=-25'd1551;
            NN[265]=25'd3413;
            NN[266]=-25'd2233;
            NN[267]=-25'd1339;
            NN[268]=-25'd5031;
            NN[269]=25'd5244;
            NN[270]=25'd11701;
            NN[271]=25'd1235;
            NN[272]=-25'd3828;
            NN[273]=-25'd4616;
            NN[274]=-25'd5306;
            NN[275]=-25'd3073;
            NN[276]=-25'd974;
            NN[277]=-25'd515;
            NN[278]=25'd61;
            NN[279]=25'd0;
            NN[280]=25'd0;
            NN[281]=25'd0;
            NN[282]=25'd473;
            NN[283]=25'd2719;
            NN[284]=25'd7359;
            NN[285]=25'd13184;
            NN[286]=25'd21869;
            NN[287]=25'd25797;
            NN[288]=25'd21605;
            NN[289]=25'd21184;
            NN[290]=25'd26759;
            NN[291]=25'd26713;
            NN[292]=25'd20918;
            NN[293]=25'd22266;
            NN[294]=25'd16434;
            NN[295]=25'd8168;
            NN[296]=25'd8764;
            NN[297]=25'd4573;
            NN[298]=-25'd4489;
            NN[299]=-25'd6175;
            NN[300]=-25'd5028;
            NN[301]=-25'd3041;
            NN[302]=-25'd2256;
            NN[303]=-25'd1044;
            NN[304]=-25'd664;
            NN[305]=-25'd120;
            NN[306]=25'd0;
            NN[307]=25'd0;
            NN[308]=25'd0;
            NN[309]=25'd0;
            NN[310]=25'd51;
            NN[311]=-25'd211;
            NN[312]=25'd704;
            NN[313]=25'd3154;
            NN[314]=25'd7136;
            NN[315]=25'd11685;
            NN[316]=25'd19533;
            NN[317]=25'd24561;
            NN[318]=25'd28160;
            NN[319]=25'd29011;
            NN[320]=25'd29480;
            NN[321]=25'd23419;
            NN[322]=25'd14392;
            NN[323]=25'd6643;
            NN[324]=25'd3956;
            NN[325]=25'd181;
            NN[326]=-25'd1292;
            NN[327]=-25'd521;
            NN[328]=-25'd2343;
            NN[329]=-25'd2866;
            NN[330]=-25'd1178;
            NN[331]=-25'd209;
            NN[332]=-25'd5;
            NN[333]=-25'd3;
            NN[334]=25'd0;
            NN[335]=25'd0;
            NN[336]=25'd0;
            NN[337]=25'd0;
            NN[338]=25'd0;
            NN[339]=25'd0;
            NN[340]=25'd9;
            NN[341]=25'd352;
            NN[342]=25'd653;
            NN[343]=25'd1294;
            NN[344]=25'd942;
            NN[345]=25'd523;
            NN[346]=25'd141;
            NN[347]=-25'd183;
            NN[348]=-25'd918;
            NN[349]=-25'd1527;
            NN[350]=-25'd2522;
            NN[351]=-25'd1955;
            NN[352]=-25'd339;
            NN[353]=-25'd548;
            NN[354]=-25'd279;
            NN[355]=-25'd578;
            NN[356]=-25'd1046;
            NN[357]=-25'd726;
            NN[358]=-25'd60;
            NN[359]=-25'd11;
            NN[360]=25'd0;
            NN[361]=25'd0;
            NN[362]=25'd0;
            NN[363]=25'd0;
            NN[364]=25'd0;
            NN[365]=25'd0;
            NN[366]=25'd0;
            NN[367]=25'd0;
            NN[368]=25'd0;
            NN[369]=25'd0;
            NN[370]=-25'd1;
            NN[371]=-25'd16;
            NN[372]=-25'd31;
            NN[373]=-25'd40;
            NN[374]=-25'd144;
            NN[375]=-25'd151;
            NN[376]=-25'd140;
            NN[377]=-25'd228;
            NN[378]=-25'd342;
            NN[379]=-25'd324;
            NN[380]=-25'd475;
            NN[381]=-25'd396;
            NN[382]=-25'd228;
            NN[383]=-25'd111;
            NN[384]=-25'd72;
            NN[385]=-25'd49;
            NN[386]=-25'd21;
            NN[387]=-25'd2;
            NN[388]=25'd0;
            NN[389]=25'd0;
            NN[390]=25'd0;
            NN[391]=25'd0;
        end
        8:begin
            NN[0]=25'd0;
            NN[1]=25'd0;
            NN[2]=25'd0;
            NN[3]=25'd0;
            NN[4]=25'd0;
            NN[5]=25'd0;
            NN[6]=25'd0;
            NN[7]=25'd0;
            NN[8]=25'd0;
            NN[9]=25'd0;
            NN[10]=25'd0;
            NN[11]=25'd0;
            NN[12]=-25'd149;
            NN[13]=-25'd329;
            NN[14]=-25'd1;
            NN[15]=25'd0;
            NN[16]=25'd0;
            NN[17]=25'd0;
            NN[18]=25'd0;
            NN[19]=25'd0;
            NN[20]=25'd0;
            NN[21]=25'd0;
            NN[22]=25'd0;
            NN[23]=25'd0;
            NN[24]=25'd0;
            NN[25]=25'd0;
            NN[26]=25'd0;
            NN[27]=25'd0;
            NN[28]=25'd0;
            NN[29]=25'd0;
            NN[30]=25'd0;
            NN[31]=25'd0;
            NN[32]=-25'd1;
            NN[33]=-25'd7;
            NN[34]=-25'd596;
            NN[35]=-25'd1403;
            NN[36]=-25'd1474;
            NN[37]=-25'd800;
            NN[38]=-25'd1606;
            NN[39]=-25'd2146;
            NN[40]=-25'd3886;
            NN[41]=-25'd2291;
            NN[42]=-25'd1236;
            NN[43]=-25'd1708;
            NN[44]=-25'd1837;
            NN[45]=-25'd922;
            NN[46]=-25'd539;
            NN[47]=-25'd285;
            NN[48]=-25'd234;
            NN[49]=-25'd519;
            NN[50]=-25'd654;
            NN[51]=-25'd193;
            NN[52]=25'd0;
            NN[53]=25'd0;
            NN[54]=25'd0;
            NN[55]=25'd0;
            NN[56]=25'd0;
            NN[57]=25'd0;
            NN[58]=25'd0;
            NN[59]=-25'd31;
            NN[60]=-25'd26;
            NN[61]=-25'd17;
            NN[62]=-25'd642;
            NN[63]=-25'd2465;
            NN[64]=-25'd3339;
            NN[65]=-25'd3922;
            NN[66]=-25'd6636;
            NN[67]=-25'd8108;
            NN[68]=-25'd10891;
            NN[69]=-25'd9630;
            NN[70]=-25'd7661;
            NN[71]=-25'd8027;
            NN[72]=-25'd8459;
            NN[73]=-25'd4918;
            NN[74]=-25'd3440;
            NN[75]=-25'd1788;
            NN[76]=-25'd1108;
            NN[77]=-25'd870;
            NN[78]=-25'd912;
            NN[79]=-25'd527;
            NN[80]=-25'd68;
            NN[81]=-25'd24;
            NN[82]=25'd0;
            NN[83]=25'd0;
            NN[84]=25'd0;
            NN[85]=25'd0;
            NN[86]=25'd0;
            NN[87]=-25'd104;
            NN[88]=-25'd72;
            NN[89]=-25'd85;
            NN[90]=-25'd1184;
            NN[91]=-25'd2853;
            NN[92]=-25'd6305;
            NN[93]=-25'd9375;
            NN[94]=-25'd10942;
            NN[95]=-25'd14233;
            NN[96]=-25'd19310;
            NN[97]=-25'd21911;
            NN[98]=-25'd18929;
            NN[99]=-25'd18528;
            NN[100]=-25'd15767;
            NN[101]=-25'd11387;
            NN[102]=-25'd7864;
            NN[103]=-25'd3398;
            NN[104]=-25'd161;
            NN[105]=25'd961;
            NN[106]=25'd594;
            NN[107]=25'd454;
            NN[108]=-25'd216;
            NN[109]=-25'd18;
            NN[110]=-25'd9;
            NN[111]=25'd0;
            NN[112]=25'd0;
            NN[113]=25'd0;
            NN[114]=-25'd2;
            NN[115]=-25'd25;
            NN[116]=25'd469;
            NN[117]=25'd532;
            NN[118]=-25'd884;
            NN[119]=-25'd3193;
            NN[120]=-25'd8098;
            NN[121]=-25'd11794;
            NN[122]=-25'd16879;
            NN[123]=-25'd19763;
            NN[124]=-25'd20773;
            NN[125]=-25'd19702;
            NN[126]=-25'd22090;
            NN[127]=-25'd20694;
            NN[128]=-25'd13439;
            NN[129]=-25'd10262;
            NN[130]=-25'd8044;
            NN[131]=-25'd602;
            NN[132]=25'd5509;
            NN[133]=25'd5889;
            NN[134]=25'd6016;
            NN[135]=25'd5730;
            NN[136]=25'd3636;
            NN[137]=25'd421;
            NN[138]=-25'd185;
            NN[139]=-25'd43;
            NN[140]=25'd0;
            NN[141]=25'd0;
            NN[142]=-25'd2;
            NN[143]=25'd42;
            NN[144]=25'd614;
            NN[145]=25'd2126;
            NN[146]=25'd2730;
            NN[147]=25'd304;
            NN[148]=-25'd2886;
            NN[149]=-25'd4330;
            NN[150]=-25'd10124;
            NN[151]=-25'd12000;
            NN[152]=-25'd14546;
            NN[153]=-25'd16754;
            NN[154]=-25'd9915;
            NN[155]=-25'd4638;
            NN[156]=25'd1114;
            NN[157]=-25'd6;
            NN[158]=25'd6610;
            NN[159]=25'd10596;
            NN[160]=25'd8523;
            NN[161]=25'd9542;
            NN[162]=25'd15479;
            NN[163]=25'd18832;
            NN[164]=25'd8111;
            NN[165]=25'd1161;
            NN[166]=-25'd395;
            NN[167]=-25'd9;
            NN[168]=25'd0;
            NN[169]=25'd0;
            NN[170]=-25'd48;
            NN[171]=-25'd403;
            NN[172]=25'd1015;
            NN[173]=25'd4559;
            NN[174]=25'd5773;
            NN[175]=25'd4929;
            NN[176]=-25'd208;
            NN[177]=-25'd963;
            NN[178]=-25'd6685;
            NN[179]=-25'd14258;
            NN[180]=-25'd17812;
            NN[181]=-25'd24501;
            NN[182]=-25'd27324;
            NN[183]=-25'd23829;
            NN[184]=-25'd19924;
            NN[185]=-25'd15863;
            NN[186]=-25'd16023;
            NN[187]=-25'd5138;
            NN[188]=-25'd3151;
            NN[189]=25'd6359;
            NN[190]=25'd23932;
            NN[191]=25'd27404;
            NN[192]=25'd12284;
            NN[193]=25'd2273;
            NN[194]=25'd890;
            NN[195]=-25'd53;
            NN[196]=25'd0;
            NN[197]=-25'd23;
            NN[198]=-25'd185;
            NN[199]=-25'd252;
            NN[200]=25'd1650;
            NN[201]=25'd6201;
            NN[202]=25'd4478;
            NN[203]=25'd3484;
            NN[204]=-25'd3067;
            NN[205]=-25'd5589;
            NN[206]=-25'd13855;
            NN[207]=-25'd20723;
            NN[208]=-25'd30859;
            NN[209]=-25'd30678;
            NN[210]=-25'd36216;
            NN[211]=-25'd39430;
            NN[212]=-25'd38677;
            NN[213]=-25'd27790;
            NN[214]=-25'd24381;
            NN[215]=-25'd17299;
            NN[216]=-25'd12467;
            NN[217]=-25'd27;
            NN[218]=25'd17444;
            NN[219]=25'd21644;
            NN[220]=25'd9408;
            NN[221]=25'd960;
            NN[222]=25'd690;
            NN[223]=-25'd53;
            NN[224]=-25'd4;
            NN[225]=-25'd305;
            NN[226]=-25'd514;
            NN[227]=-25'd1032;
            NN[228]=25'd264;
            NN[229]=25'd4789;
            NN[230]=25'd1266;
            NN[231]=-25'd3002;
            NN[232]=-25'd10246;
            NN[233]=-25'd3942;
            NN[234]=-25'd14389;
            NN[235]=-25'd15078;
            NN[236]=-25'd23362;
            NN[237]=-25'd23559;
            NN[238]=-25'd38538;
            NN[239]=-25'd41124;
            NN[240]=-25'd34093;
            NN[241]=-25'd20865;
            NN[242]=-25'd13775;
            NN[243]=-25'd10457;
            NN[244]=-25'd7792;
            NN[245]=-25'd3241;
            NN[246]=25'd4777;
            NN[247]=25'd7047;
            NN[248]=25'd1080;
            NN[249]=-25'd2594;
            NN[250]=-25'd2092;
            NN[251]=-25'd83;
            NN[252]=-25'd29;
            NN[253]=-25'd356;
            NN[254]=-25'd858;
            NN[255]=-25'd3695;
            NN[256]=-25'd4297;
            NN[257]=-25'd1215;
            NN[258]=-25'd7018;
            NN[259]=-25'd8569;
            NN[260]=-25'd6844;
            NN[261]=-25'd1989;
            NN[262]=-25'd9966;
            NN[263]=-25'd8441;
            NN[264]=-25'd7322;
            NN[265]=-25'd14071;
            NN[266]=-25'd48308;
            NN[267]=-25'd39744;
            NN[268]=-25'd11983;
            NN[269]=-25'd3747;
            NN[270]=-25'd4520;
            NN[271]=-25'd4392;
            NN[272]=-25'd3856;
            NN[273]=-25'd3738;
            NN[274]=-25'd3528;
            NN[275]=-25'd7952;
            NN[276]=-25'd14162;
            NN[277]=-25'd9392;
            NN[278]=-25'd2914;
            NN[279]=-25'd256;
            NN[280]=-25'd34;
            NN[281]=-25'd329;
            NN[282]=-25'd1411;
            NN[283]=-25'd4039;
            NN[284]=-25'd5077;
            NN[285]=-25'd5604;
            NN[286]=-25'd10595;
            NN[287]=-25'd7064;
            NN[288]=-25'd336;
            NN[289]=25'd9952;
            NN[290]=25'd5133;
            NN[291]=25'd5171;
            NN[292]=25'd11797;
            NN[293]=-25'd18250;
            NN[294]=-25'd53332;
            NN[295]=-25'd22647;
            NN[296]=25'd2337;
            NN[297]=25'd7661;
            NN[298]=-25'd3190;
            NN[299]=-25'd1212;
            NN[300]=-25'd10239;
            NN[301]=-25'd9159;
            NN[302]=-25'd12309;
            NN[303]=-25'd19696;
            NN[304]=-25'd15898;
            NN[305]=-25'd9559;
            NN[306]=-25'd2658;
            NN[307]=-25'd55;
            NN[308]=-25'd5;
            NN[309]=-25'd675;
            NN[310]=-25'd3320;
            NN[311]=-25'd4231;
            NN[312]=-25'd7509;
            NN[313]=-25'd6773;
            NN[314]=-25'd4147;
            NN[315]=25'd1541;
            NN[316]=25'd13891;
            NN[317]=25'd20573;
            NN[318]=25'd24307;
            NN[319]=25'd25197;
            NN[320]=25'd24352;
            NN[321]=-25'd30680;
            NN[322]=-25'd47241;
            NN[323]=-25'd2456;
            NN[324]=25'd26744;
            NN[325]=25'd11743;
            NN[326]=-25'd3229;
            NN[327]=-25'd6367;
            NN[328]=-25'd12233;
            NN[329]=-25'd12370;
            NN[330]=-25'd14836;
            NN[331]=-25'd17010;
            NN[332]=-25'd12197;
            NN[333]=-25'd4901;
            NN[334]=-25'd630;
            NN[335]=-25'd32;
            NN[336]=-25'd2;
            NN[337]=-25'd956;
            NN[338]=-25'd3592;
            NN[339]=-25'd5702;
            NN[340]=-25'd9405;
            NN[341]=-25'd4732;
            NN[342]=25'd7685;
            NN[343]=25'd18237;
            NN[344]=25'd26610;
            NN[345]=25'd25877;
            NN[346]=25'd38101;
            NN[347]=25'd48438;
            NN[348]=25'd40573;
            NN[349]=-25'd10227;
            NN[350]=-25'd27444;
            NN[351]=25'd11953;
            NN[352]=25'd30507;
            NN[353]=25'd14118;
            NN[354]=25'd3535;
            NN[355]=25'd1128;
            NN[356]=-25'd695;
            NN[357]=-25'd561;
            NN[358]=-25'd4488;
            NN[359]=-25'd9077;
            NN[360]=-25'd4712;
            NN[361]=-25'd1314;
            NN[362]=-25'd570;
            NN[363]=-25'd196;
            NN[364]=25'd0;
            NN[365]=-25'd731;
            NN[366]=-25'd2103;
            NN[367]=-25'd4285;
            NN[368]=-25'd3799;
            NN[369]=25'd7767;
            NN[370]=25'd24599;
            NN[371]=25'd28656;
            NN[372]=25'd30401;
            NN[373]=25'd31522;
            NN[374]=25'd42520;
            NN[375]=25'd52938;
            NN[376]=25'd30433;
            NN[377]=-25'd6976;
            NN[378]=-25'd10720;
            NN[379]=25'd15730;
            NN[380]=25'd27004;
            NN[381]=25'd26159;
            NN[382]=25'd15486;
            NN[383]=25'd10685;
            NN[384]=25'd14303;
            NN[385]=25'd6777;
            NN[386]=25'd2562;
            NN[387]=-25'd1937;
            NN[388]=-25'd3905;
            NN[389]=-25'd157;
            NN[390]=-25'd393;
            NN[391]=-25'd609;
        end
        9:begin
            NN[0]=-25'd2;
            NN[1]=-25'd402;
            NN[2]=-25'd926;
            NN[3]=-25'd703;
            NN[4]=25'd8573;
            NN[5]=25'd20759;
            NN[6]=25'd29274;
            NN[7]=25'd33470;
            NN[8]=25'd29851;
            NN[9]=25'd27713;
            NN[10]=25'd35412;
            NN[11]=25'd37767;
            NN[12]=25'd19314;
            NN[13]=-25'd6755;
            NN[14]=-25'd5371;
            NN[15]=25'd12620;
            NN[16]=25'd34450;
            NN[17]=25'd40142;
            NN[18]=25'd25670;
            NN[19]=25'd25988;
            NN[20]=25'd18094;
            NN[21]=25'd6603;
            NN[22]=25'd3262;
            NN[23]=-25'd1459;
            NN[24]=-25'd4439;
            NN[25]=-25'd1682;
            NN[26]=-25'd986;
            NN[27]=-25'd70;
            NN[28]=-25'd1;
            NN[29]=-25'd19;
            NN[30]=25'd162;
            NN[31]=25'd1292;
            NN[32]=25'd8263;
            NN[33]=25'd16908;
            NN[34]=25'd23979;
            NN[35]=25'd30701;
            NN[36]=25'd33445;
            NN[37]=25'd27916;
            NN[38]=25'd21492;
            NN[39]=25'd22820;
            NN[40]=25'd10928;
            NN[41]=-25'd5519;
            NN[42]=25'd3336;
            NN[43]=25'd25228;
            NN[44]=25'd44134;
            NN[45]=25'd36959;
            NN[46]=25'd20177;
            NN[47]=25'd18755;
            NN[48]=25'd5123;
            NN[49]=25'd178;
            NN[50]=25'd1216;
            NN[51]=-25'd4638;
            NN[52]=-25'd10395;
            NN[53]=-25'd4775;
            NN[54]=25'd330;
            NN[55]=-25'd107;
            NN[56]=-25'd1;
            NN[57]=-25'd9;
            NN[58]=-25'd455;
            NN[59]=-25'd2440;
            NN[60]=-25'd2391;
            NN[61]=25'd5845;
            NN[62]=25'd14287;
            NN[63]=25'd27853;
            NN[64]=25'd30956;
            NN[65]=25'd22110;
            NN[66]=25'd3439;
            NN[67]=-25'd404;
            NN[68]=25'd5263;
            NN[69]=25'd6102;
            NN[70]=25'd23458;
            NN[71]=25'd43946;
            NN[72]=25'd39988;
            NN[73]=25'd25061;
            NN[74]=25'd16923;
            NN[75]=25'd8422;
            NN[76]=25'd7819;
            NN[77]=25'd2813;
            NN[78]=-25'd6061;
            NN[79]=-25'd9218;
            NN[80]=-25'd9394;
            NN[81]=-25'd5502;
            NN[82]=-25'd1671;
            NN[83]=-25'd64;
            NN[84]=25'd0;
            NN[85]=-25'd3;
            NN[86]=-25'd547;
            NN[87]=-25'd5727;
            NN[88]=-25'd5548;
            NN[89]=-25'd3968;
            NN[90]=25'd2518;
            NN[91]=25'd14652;
            NN[92]=25'd20141;
            NN[93]=25'd12621;
            NN[94]=25'd2631;
            NN[95]=-25'd1356;
            NN[96]=25'd7105;
            NN[97]=25'd21737;
            NN[98]=25'd39780;
            NN[99]=25'd40453;
            NN[100]=25'd27367;
            NN[101]=25'd13730;
            NN[102]=25'd10407;
            NN[103]=-25'd3186;
            NN[104]=-25'd1619;
            NN[105]=-25'd3151;
            NN[106]=-25'd11432;
            NN[107]=-25'd9696;
            NN[108]=-25'd8198;
            NN[109]=-25'd6177;
            NN[110]=-25'd926;
            NN[111]=-25'd315;
            NN[112]=-25'd72;
            NN[113]=25'd0;
            NN[114]=-25'd462;
            NN[115]=-25'd5053;
            NN[116]=-25'd6779;
            NN[117]=-25'd7524;
            NN[118]=-25'd9217;
            NN[119]=-25'd4139;
            NN[120]=-25'd557;
            NN[121]=-25'd4554;
            NN[122]=-25'd16530;
            NN[123]=-25'd12878;
            NN[124]=25'd3132;
            NN[125]=25'd15713;
            NN[126]=25'd24746;
            NN[127]=25'd21527;
            NN[128]=25'd13831;
            NN[129]=-25'd7163;
            NN[130]=-25'd5685;
            NN[131]=-25'd11341;
            NN[132]=-25'd8935;
            NN[133]=-25'd10505;
            NN[134]=-25'd17991;
            NN[135]=-25'd12217;
            NN[136]=-25'd8237;
            NN[137]=-25'd5831;
            NN[138]=-25'd440;
            NN[139]=-25'd1;
            NN[140]=25'd0;
            NN[141]=-25'd80;
            NN[142]=-25'd561;
            NN[143]=-25'd2356;
            NN[144]=-25'd6931;
            NN[145]=-25'd8225;
            NN[146]=-25'd15728;
            NN[147]=-25'd20792;
            NN[148]=-25'd25768;
            NN[149]=-25'd31381;
            NN[150]=-25'd34907;
            NN[151]=-25'd27800;
            NN[152]=-25'd27239;
            NN[153]=-25'd11954;
            NN[154]=25'd5942;
            NN[155]=25'd4717;
            NN[156]=-25'd2299;
            NN[157]=-25'd10183;
            NN[158]=-25'd12092;
            NN[159]=-25'd14766;
            NN[160]=-25'd12793;
            NN[161]=-25'd11328;
            NN[162]=-25'd18863;
            NN[163]=-25'd12274;
            NN[164]=-25'd7549;
            NN[165]=-25'd2614;
            NN[166]=-25'd86;
            NN[167]=25'd0;
            NN[168]=25'd0;
            NN[169]=-25'd3;
            NN[170]=-25'd341;
            NN[171]=-25'd2778;
            NN[172]=-25'd6614;
            NN[173]=-25'd12001;
            NN[174]=-25'd19919;
            NN[175]=-25'd29920;
            NN[176]=-25'd37241;
            NN[177]=-25'd38133;
            NN[178]=-25'd34985;
            NN[179]=-25'd25090;
            NN[180]=-25'd23008;
            NN[181]=-25'd20851;
            NN[182]=-25'd7663;
            NN[183]=-25'd1065;
            NN[184]=-25'd2793;
            NN[185]=-25'd6342;
            NN[186]=-25'd10293;
            NN[187]=-25'd9859;
            NN[188]=-25'd8206;
            NN[189]=-25'd7478;
            NN[190]=-25'd12327;
            NN[191]=-25'd9426;
            NN[192]=-25'd4223;
            NN[193]=-25'd1861;
            NN[194]=-25'd44;
            NN[195]=25'd0;
            NN[196]=25'd0;
            NN[197]=25'd0;
            NN[198]=-25'd71;
            NN[199]=-25'd1881;
            NN[200]=-25'd4272;
            NN[201]=-25'd8380;
            NN[202]=-25'd17883;
            NN[203]=-25'd24932;
            NN[204]=-25'd22582;
            NN[205]=-25'd23155;
            NN[206]=-25'd23041;
            NN[207]=-25'd14238;
            NN[208]=-25'd13095;
            NN[209]=-25'd15705;
            NN[210]=-25'd7860;
            NN[211]=25'd1276;
            NN[212]=-25'd4757;
            NN[213]=-25'd1574;
            NN[214]=-25'd4320;
            NN[215]=25'd2549;
            NN[216]=25'd1263;
            NN[217]=-25'd1440;
            NN[218]=-25'd4906;
            NN[219]=-25'd3742;
            NN[220]=-25'd2552;
            NN[221]=-25'd1543;
            NN[222]=-25'd64;
            NN[223]=25'd0;
            NN[224]=25'd0;
            NN[225]=25'd0;
            NN[226]=-25'd33;
            NN[227]=-25'd1319;
            NN[228]=-25'd2739;
            NN[229]=-25'd6052;
            NN[230]=-25'd11168;
            NN[231]=-25'd15874;
            NN[232]=-25'd15306;
            NN[233]=-25'd16618;
            NN[234]=-25'd12241;
            NN[235]=-25'd9460;
            NN[236]=-25'd9947;
            NN[237]=-25'd9325;
            NN[238]=-25'd8346;
            NN[239]=-25'd2447;
            NN[240]=-25'd3697;
            NN[241]=25'd2938;
            NN[242]=25'd6555;
            NN[243]=25'd16537;
            NN[244]=25'd10528;
            NN[245]=25'd9069;
            NN[246]=25'd923;
            NN[247]=-25'd2695;
            NN[248]=-25'd1810;
            NN[249]=-25'd1049;
            NN[250]=25'd20;
            NN[251]=25'd0;
            NN[252]=25'd0;
            NN[253]=25'd0;
            NN[254]=-25'd10;
            NN[255]=-25'd412;
            NN[256]=-25'd1537;
            NN[257]=-25'd3779;
            NN[258]=-25'd5441;
            NN[259]=-25'd7375;
            NN[260]=-25'd7748;
            NN[261]=-25'd7591;
            NN[262]=-25'd5753;
            NN[263]=-25'd2817;
            NN[264]=-25'd9034;
            NN[265]=-25'd6699;
            NN[266]=-25'd3486;
            NN[267]=-25'd856;
            NN[268]=25'd2420;
            NN[269]=25'd6548;
            NN[270]=25'd15534;
            NN[271]=25'd16898;
            NN[272]=25'd15043;
            NN[273]=25'd9415;
            NN[274]=25'd220;
            NN[275]=-25'd1924;
            NN[276]=-25'd1614;
            NN[277]=-25'd258;
            NN[278]=25'd26;
            NN[279]=25'd0;
            NN[280]=25'd0;
            NN[281]=25'd0;
            NN[282]=25'd0;
            NN[283]=-25'd25;
            NN[284]=-25'd877;
            NN[285]=-25'd1604;
            NN[286]=-25'd3104;
            NN[287]=-25'd3582;
            NN[288]=-25'd4373;
            NN[289]=-25'd3552;
            NN[290]=-25'd2610;
            NN[291]=-25'd1044;
            NN[292]=-25'd9660;
            NN[293]=-25'd10691;
            NN[294]=-25'd7407;
            NN[295]=-25'd7893;
            NN[296]=-25'd3474;
            NN[297]=-25'd3787;
            NN[298]=25'd2627;
            NN[299]=25'd7243;
            NN[300]=25'd5240;
            NN[301]=25'd2607;
            NN[302]=-25'd255;
            NN[303]=-25'd1139;
            NN[304]=-25'd983;
            NN[305]=-25'd22;
            NN[306]=-25'd2;
            NN[307]=25'd0;
            NN[308]=25'd0;
            NN[309]=25'd0;
            NN[310]=-25'd1;
            NN[311]=-25'd3;
            NN[312]=-25'd295;
            NN[313]=-25'd1848;
            NN[314]=-25'd3571;
            NN[315]=-25'd7111;
            NN[316]=-25'd13260;
            NN[317]=-25'd13994;
            NN[318]=-25'd12588;
            NN[319]=-25'd18583;
            NN[320]=-25'd25330;
            NN[321]=-25'd21247;
            NN[322]=-25'd20379;
            NN[323]=-25'd22146;
            NN[324]=-25'd24409;
            NN[325]=-25'd24765;
            NN[326]=-25'd20247;
            NN[327]=-25'd16052;
            NN[328]=-25'd9440;
            NN[329]=-25'd4917;
            NN[330]=-25'd2038;
            NN[331]=-25'd1128;
            NN[332]=-25'd724;
            NN[333]=-25'd109;
            NN[334]=-25'd2;
            NN[335]=25'd0;
            NN[336]=25'd0;
            NN[337]=25'd0;
            NN[338]=25'd0;
            NN[339]=25'd0;
            NN[340]=-25'd155;
            NN[341]=-25'd618;
            NN[342]=-25'd1642;
            NN[343]=-25'd3436;
            NN[344]=-25'd6152;
            NN[345]=-25'd10071;
            NN[346]=-25'd11598;
            NN[347]=-25'd14752;
            NN[348]=-25'd17616;
            NN[349]=-25'd17882;
            NN[350]=-25'd20503;
            NN[351]=-25'd18763;
            NN[352]=-25'd17315;
            NN[353]=-25'd14410;
            NN[354]=-25'd13629;
            NN[355]=-25'd9875;
            NN[356]=-25'd4770;
            NN[357]=-25'd2253;
            NN[358]=-25'd1063;
            NN[359]=-25'd38;
            NN[360]=-25'd19;
            NN[361]=25'd0;
            NN[362]=25'd0;
            NN[363]=25'd0;
            NN[364]=25'd0;
            NN[365]=25'd0;
            NN[366]=25'd0;
            NN[367]=25'd0;
            NN[368]=25'd0;
            NN[369]=25'd0;
            NN[370]=-25'd70;
            NN[371]=-25'd436;
            NN[372]=-25'd595;
            NN[373]=-25'd499;
            NN[374]=-25'd967;
            NN[375]=-25'd847;
            NN[376]=-25'd1181;
            NN[377]=-25'd1016;
            NN[378]=-25'd1969;
            NN[379]=-25'd1167;
            NN[380]=-25'd1426;
            NN[381]=-25'd1222;
            NN[382]=-25'd1222;
            NN[383]=-25'd766;
            NN[384]=-25'd162;
            NN[385]=-25'd79;
            NN[386]=-25'd109;
            NN[387]=-25'd23;
            NN[388]=25'd0;
            NN[389]=25'd0;
            NN[390]=25'd0;
            NN[391]=25'd0;
        end
        10:begin
            NN[0]=25'd0;
            NN[1]=25'd0;
            NN[2]=25'd0;
            NN[3]=25'd0;
            NN[4]=25'd0;
            NN[5]=25'd0;
            NN[6]=25'd0;
            NN[7]=25'd0;
            NN[8]=25'd0;
            NN[9]=25'd0;
            NN[10]=25'd0;
            NN[11]=25'd0;
            NN[12]=-25'd3;
            NN[13]=-25'd7;
            NN[14]=25'd0;
            NN[15]=25'd0;
            NN[16]=25'd0;
            NN[17]=25'd0;
            NN[18]=25'd0;
            NN[19]=25'd0;
            NN[20]=25'd0;
            NN[21]=25'd0;
            NN[22]=25'd0;
            NN[23]=25'd0;
            NN[24]=25'd0;
            NN[25]=25'd0;
            NN[26]=25'd0;
            NN[27]=25'd0;
            NN[28]=25'd0;
            NN[29]=25'd0;
            NN[30]=25'd0;
            NN[31]=25'd0;
            NN[32]=25'd0;
            NN[33]=25'd0;
            NN[34]=25'd0;
            NN[35]=-25'd1;
            NN[36]=-25'd2;
            NN[37]=-25'd38;
            NN[38]=-25'd105;
            NN[39]=-25'd36;
            NN[40]=-25'd121;
            NN[41]=-25'd122;
            NN[42]=-25'd69;
            NN[43]=-25'd76;
            NN[44]=-25'd122;
            NN[45]=-25'd62;
            NN[46]=-25'd70;
            NN[47]=-25'd58;
            NN[48]=-25'd29;
            NN[49]=-25'd8;
            NN[50]=25'd0;
            NN[51]=25'd0;
            NN[52]=25'd0;
            NN[53]=25'd0;
            NN[54]=25'd0;
            NN[55]=25'd0;
            NN[56]=25'd0;
            NN[57]=25'd0;
            NN[58]=25'd0;
            NN[59]=-25'd2;
            NN[60]=25'd0;
            NN[61]=25'd0;
            NN[62]=-25'd2;
            NN[63]=-25'd77;
            NN[64]=-25'd105;
            NN[65]=-25'd421;
            NN[66]=-25'd983;
            NN[67]=-25'd1769;
            NN[68]=-25'd2004;
            NN[69]=-25'd2334;
            NN[70]=-25'd2816;
            NN[71]=-25'd2224;
            NN[72]=-25'd940;
            NN[73]=25'd116;
            NN[74]=-25'd64;
            NN[75]=-25'd507;
            NN[76]=-25'd1323;
            NN[77]=-25'd1494;
            NN[78]=-25'd906;
            NN[79]=-25'd567;
            NN[80]=-25'd223;
            NN[81]=-25'd37;
            NN[82]=25'd0;
            NN[83]=25'd0;
            NN[84]=25'd0;
            NN[85]=25'd0;
            NN[86]=25'd0;
            NN[87]=-25'd4;
            NN[88]=25'd202;
            NN[89]=-25'd378;
            NN[90]=-25'd390;
            NN[91]=-25'd1157;
            NN[92]=-25'd1519;
            NN[93]=-25'd2534;
            NN[94]=-25'd2514;
            NN[95]=-25'd4741;
            NN[96]=-25'd4764;
            NN[97]=-25'd5903;
            NN[98]=-25'd5163;
            NN[99]=-25'd985;
            NN[100]=25'd425;
            NN[101]=25'd4709;
            NN[102]=25'd7253;
            NN[103]=25'd5338;
            NN[104]=25'd4730;
            NN[105]=25'd3674;
            NN[106]=25'd1813;
            NN[107]=-25'd1853;
            NN[108]=-25'd1556;
            NN[109]=25'd471;
            NN[110]=25'd103;
            NN[111]=25'd0;
            NN[112]=25'd0;
            NN[113]=25'd0;
            NN[114]=-25'd23;
            NN[115]=-25'd163;
            NN[116]=-25'd1067;
            NN[117]=-25'd3832;
            NN[118]=-25'd5603;
            NN[119]=-25'd7241;
            NN[120]=-25'd12434;
            NN[121]=-25'd12513;
            NN[122]=-25'd8613;
            NN[123]=-25'd6161;
            NN[124]=-25'd10248;
            NN[125]=-25'd15454;
            NN[126]=-25'd6720;
            NN[127]=25'd7561;
            NN[128]=25'd9746;
            NN[129]=25'd12105;
            NN[130]=25'd11690;
            NN[131]=25'd3367;
            NN[132]=-25'd1930;
            NN[133]=25'd8696;
            NN[134]=25'd9556;
            NN[135]=25'd11105;
            NN[136]=25'd8390;
            NN[137]=25'd2759;
            NN[138]=25'd478;
            NN[139]=-25'd62;
            NN[140]=25'd0;
            NN[141]=25'd0;
            NN[142]=-25'd125;
            NN[143]=-25'd967;
            NN[144]=-25'd3950;
            NN[145]=-25'd7881;
            NN[146]=-25'd11134;
            NN[147]=-25'd10098;
            NN[148]=-25'd8709;
            NN[149]=-25'd1926;
            NN[150]=25'd2297;
            NN[151]=25'd3209;
            NN[152]=-25'd3079;
            NN[153]=-25'd5787;
            NN[154]=-25'd6291;
            NN[155]=-25'd6856;
            NN[156]=25'd1237;
            NN[157]=25'd6664;
            NN[158]=25'd7394;
            NN[159]=25'd3197;
            NN[160]=25'd9640;
            NN[161]=25'd11411;
            NN[162]=25'd19447;
            NN[163]=25'd23611;
            NN[164]=25'd18534;
            NN[165]=25'd9410;
            NN[166]=25'd2095;
            NN[167]=25'd169;
            NN[168]=25'd0;
            NN[169]=25'd0;
            NN[170]=25'd20;
            NN[171]=-25'd2836;
            NN[172]=-25'd7136;
            NN[173]=-25'd10153;
            NN[174]=-25'd10970;
            NN[175]=-25'd4753;
            NN[176]=25'd578;
            NN[177]=25'd4229;
            NN[178]=25'd7222;
            NN[179]=25'd3984;
            NN[180]=25'd493;
            NN[181]=-25'd1786;
            NN[182]=25'd3415;
            NN[183]=-25'd4924;
            NN[184]=-25'd6529;
            NN[185]=-25'd2480;
            NN[186]=25'd5246;
            NN[187]=25'd11528;
            NN[188]=25'd11173;
            NN[189]=25'd8606;
            NN[190]=25'd19088;
            NN[191]=25'd31867;
            NN[192]=25'd35876;
            NN[193]=25'd20830;
            NN[194]=25'd6429;
            NN[195]=25'd1023;
            NN[196]=25'd0;
            NN[197]=-25'd24;
            NN[198]=-25'd592;
            NN[199]=-25'd3776;
            NN[200]=-25'd13576;
            NN[201]=-25'd15346;
            NN[202]=-25'd11388;
            NN[203]=-25'd1968;
            NN[204]=25'd8131;
            NN[205]=25'd10402;
            NN[206]=25'd12053;
            NN[207]=25'd11192;
            NN[208]=25'd4491;
            NN[209]=-25'd5484;
            NN[210]=25'd2967;
            NN[211]=-25'd9174;
            NN[212]=-25'd1201;
            NN[213]=25'd4982;
            NN[214]=25'd7639;
            NN[215]=25'd9728;
            NN[216]=25'd9997;
            NN[217]=25'd9124;
            NN[218]=25'd16882;
            NN[219]=25'd36600;
            NN[220]=25'd47116;
            NN[221]=25'd34254;
            NN[222]=25'd8057;
            NN[223]=25'd794;
            NN[224]=25'd0;
            NN[225]=-25'd53;
            NN[226]=-25'd787;
            NN[227]=-25'd4545;
            NN[228]=-25'd17973;
            NN[229]=-25'd17228;
            NN[230]=-25'd11915;
            NN[231]=-25'd5147;
            NN[232]=25'd9800;
            NN[233]=25'd8830;
            NN[234]=25'd8486;
            NN[235]=25'd11691;
            NN[236]=-25'd238;
            NN[237]=-25'd9575;
            NN[238]=-25'd11828;
            NN[239]=-25'd19902;
            NN[240]=-25'd11737;
            NN[241]=-25'd4646;
            NN[242]=-25'd2828;
            NN[243]=25'd2560;
            NN[244]=25'd10790;
            NN[245]=25'd13274;
            NN[246]=25'd18903;
            NN[247]=25'd48266;
            NN[248]=25'd64587;
            NN[249]=25'd42820;
            NN[250]=25'd11052;
            NN[251]=25'd727;
            NN[252]=-25'd2;
            NN[253]=-25'd57;
            NN[254]=-25'd479;
            NN[255]=-25'd4979;
            NN[256]=-25'd15364;
            NN[257]=-25'd15708;
            NN[258]=-25'd8248;
            NN[259]=25'd4709;
            NN[260]=25'd15483;
            NN[261]=25'd15309;
            NN[262]=25'd18258;
            NN[263]=25'd25976;
            NN[264]=25'd10181;
            NN[265]=-25'd4226;
            NN[266]=-25'd18135;
            NN[267]=-25'd26505;
            NN[268]=-25'd26313;
            NN[269]=-25'd19337;
            NN[270]=-25'd13188;
            NN[271]=-25'd6027;
            NN[272]=25'd5258;
            NN[273]=25'd19844;
            NN[274]=25'd27704;
            NN[275]=25'd53164;
            NN[276]=25'd75405;
            NN[277]=25'd49915;
            NN[278]=25'd11336;
            NN[279]=25'd770;
            NN[280]=-25'd2;
            NN[281]=-25'd56;
            NN[282]=-25'd440;
            NN[283]=-25'd4183;
            NN[284]=-25'd7931;
            NN[285]=-25'd7660;
            NN[286]=25'd985;
            NN[287]=25'd13815;
            NN[288]=25'd22950;
            NN[289]=25'd28425;
            NN[290]=25'd26406;
            NN[291]=25'd25948;
            NN[292]=25'd22081;
            NN[293]=25'd13651;
            NN[294]=25'd1393;
            NN[295]=-25'd10190;
            NN[296]=-25'd17053;
            NN[297]=-25'd24752;
            NN[298]=-25'd24174;
            NN[299]=-25'd20000;
            NN[300]=-25'd8978;
            NN[301]=25'd426;
            NN[302]=25'd8136;
            NN[303]=25'd32232;
            NN[304]=25'd57622;
            NN[305]=25'd46359;
            NN[306]=25'd11887;
            NN[307]=25'd328;
            NN[308]=-25'd3;
            NN[309]=-25'd272;
            NN[310]=-25'd755;
            NN[311]=-25'd4187;
            NN[312]=-25'd3251;
            NN[313]=25'd737;
            NN[314]=25'd12417;
            NN[315]=25'd15600;
            NN[316]=25'd15310;
            NN[317]=25'd17616;
            NN[318]=25'd17734;
            NN[319]=25'd18875;
            NN[320]=25'd29380;
            NN[321]=25'd34431;
            NN[322]=25'd13896;
            NN[323]=-25'd5169;
            NN[324]=-25'd13034;
            NN[325]=-25'd19916;
            NN[326]=-25'd22257;
            NN[327]=-25'd34300;
            NN[328]=-25'd42179;
            NN[329]=-25'd35495;
            NN[330]=-25'd32171;
            NN[331]=-25'd11253;
            NN[332]=25'd11229;
            NN[333]=25'd21035;
            NN[334]=25'd6044;
            NN[335]=25'd196;
            NN[336]=-25'd2;
            NN[337]=-25'd331;
            NN[338]=-25'd645;
            NN[339]=-25'd1653;
            NN[340]=25'd16;
            NN[341]=25'd5919;
            NN[342]=25'd13740;
            NN[343]=25'd14245;
            NN[344]=25'd10234;
            NN[345]=25'd4460;
            NN[346]=25'd19143;
            NN[347]=25'd26936;
            NN[348]=25'd32223;
            NN[349]=25'd31030;
            NN[350]=25'd4950;
            NN[351]=-25'd11205;
            NN[352]=-25'd28129;
            NN[353]=-25'd28774;
            NN[354]=-25'd26120;
            NN[355]=-25'd30445;
            NN[356]=-25'd38755;
            NN[357]=-25'd50558;
            NN[358]=-25'd54652;
            NN[359]=-25'd41908;
            NN[360]=-25'd24245;
            NN[361]=25'd247;
            NN[362]=25'd2206;
            NN[363]=-25'd58;
            NN[364]=25'd0;
            NN[365]=-25'd79;
            NN[366]=-25'd241;
            NN[367]=25'd16;
            NN[368]=25'd2404;
            NN[369]=25'd9513;
            NN[370]=25'd7208;
            NN[371]=25'd13729;
            NN[372]=25'd10877;
            NN[373]=25'd12427;
            NN[374]=25'd23251;
            NN[375]=25'd27085;
            NN[376]=25'd30833;
            NN[377]=25'd20980;
            NN[378]=25'd1329;
            NN[379]=-25'd20863;
            NN[380]=-25'd32439;
            NN[381]=-25'd21074;
            NN[382]=-25'd12795;
            NN[383]=-25'd12083;
            NN[384]=-25'd14013;
            NN[385]=-25'd27039;
            NN[386]=-25'd32231;
            NN[387]=-25'd35206;
            NN[388]=-25'd22634;
            NN[389]=-25'd3571;
            NN[390]=-25'd233;
            NN[391]=-25'd442;
        end
        11:begin
            NN[0]=25'd175;
            NN[1]=-25'd50;
            NN[2]=-25'd109;
            NN[3]=25'd212;
            NN[4]=25'd1717;
            NN[5]=25'd2510;
            NN[6]=-25'd327;
            NN[7]=25'd2227;
            NN[8]=25'd7958;
            NN[9]=25'd21580;
            NN[10]=25'd26942;
            NN[11]=25'd14953;
            NN[12]=25'd12605;
            NN[13]=25'd6587;
            NN[14]=-25'd7691;
            NN[15]=-25'd18710;
            NN[16]=-25'd25721;
            NN[17]=-25'd20527;
            NN[18]=-25'd11432;
            NN[19]=-25'd11869;
            NN[20]=-25'd5993;
            NN[21]=-25'd10788;
            NN[22]=-25'd11216;
            NN[23]=-25'd16690;
            NN[24]=-25'd14294;
            NN[25]=-25'd4667;
            NN[26]=-25'd690;
            NN[27]=-25'd32;
            NN[28]=25'd55;
            NN[29]=-25'd56;
            NN[30]=-25'd123;
            NN[31]=-25'd473;
            NN[32]=-25'd1282;
            NN[33]=-25'd7325;
            NN[34]=-25'd9689;
            NN[35]=-25'd13746;
            NN[36]=-25'd1614;
            NN[37]=25'd14206;
            NN[38]=25'd15594;
            NN[39]=25'd13137;
            NN[40]=25'd12978;
            NN[41]=-25'd896;
            NN[42]=-25'd20763;
            NN[43]=-25'd22021;
            NN[44]=-25'd22009;
            NN[45]=-25'd17998;
            NN[46]=-25'd759;
            NN[47]=-25'd8543;
            NN[48]=-25'd7160;
            NN[49]=-25'd4016;
            NN[50]=-25'd4940;
            NN[51]=-25'd4528;
            NN[52]=-25'd5824;
            NN[53]=-25'd3567;
            NN[54]=-25'd1015;
            NN[55]=-25'd283;
            NN[56]=-25'd13;
            NN[57]=-25'd28;
            NN[58]=-25'd269;
            NN[59]=25'd216;
            NN[60]=-25'd1812;
            NN[61]=-25'd7874;
            NN[62]=-25'd11733;
            NN[63]=-25'd24671;
            NN[64]=-25'd24317;
            NN[65]=-25'd19875;
            NN[66]=-25'd11939;
            NN[67]=-25'd9989;
            NN[68]=-25'd4108;
            NN[69]=-25'd12380;
            NN[70]=-25'd21697;
            NN[71]=-25'd14341;
            NN[72]=-25'd15928;
            NN[73]=-25'd8659;
            NN[74]=-25'd3294;
            NN[75]=-25'd1088;
            NN[76]=25'd781;
            NN[77]=-25'd1790;
            NN[78]=25'd1663;
            NN[79]=25'd1837;
            NN[80]=-25'd729;
            NN[81]=-25'd3297;
            NN[82]=-25'd1226;
            NN[83]=-25'd407;
            NN[84]=25'd0;
            NN[85]=-25'd14;
            NN[86]=-25'd455;
            NN[87]=25'd683;
            NN[88]=25'd1421;
            NN[89]=25'd7220;
            NN[90]=25'd15745;
            NN[91]=-25'd9524;
            NN[92]=-25'd23033;
            NN[93]=-25'd24331;
            NN[94]=-25'd28171;
            NN[95]=-25'd24275;
            NN[96]=-25'd27087;
            NN[97]=-25'd25814;
            NN[98]=-25'd18427;
            NN[99]=-25'd9432;
            NN[100]=-25'd2358;
            NN[101]=25'd3745;
            NN[102]=25'd8761;
            NN[103]=25'd5865;
            NN[104]=25'd7956;
            NN[105]=25'd3502;
            NN[106]=-25'd1794;
            NN[107]=25'd4399;
            NN[108]=25'd3920;
            NN[109]=-25'd3387;
            NN[110]=-25'd717;
            NN[111]=-25'd83;
            NN[112]=-25'd10;
            NN[113]=-25'd4;
            NN[114]=-25'd409;
            NN[115]=25'd617;
            NN[116]=25'd6721;
            NN[117]=25'd16085;
            NN[118]=25'd34013;
            NN[119]=25'd15187;
            NN[120]=25'd708;
            NN[121]=-25'd10735;
            NN[122]=-25'd17637;
            NN[123]=-25'd14472;
            NN[124]=-25'd9384;
            NN[125]=-25'd5368;
            NN[126]=25'd215;
            NN[127]=25'd605;
            NN[128]=25'd1158;
            NN[129]=25'd5826;
            NN[130]=25'd1458;
            NN[131]=25'd6476;
            NN[132]=25'd11278;
            NN[133]=25'd4599;
            NN[134]=25'd2225;
            NN[135]=25'd6546;
            NN[136]=25'd7186;
            NN[137]=-25'd1950;
            NN[138]=-25'd419;
            NN[139]=-25'd194;
            NN[140]=25'd0;
            NN[141]=-25'd18;
            NN[142]=-25'd525;
            NN[143]=-25'd639;
            NN[144]=25'd7444;
            NN[145]=25'd19580;
            NN[146]=25'd29191;
            NN[147]=25'd18166;
            NN[148]=25'd19982;
            NN[149]=25'd10139;
            NN[150]=25'd2570;
            NN[151]=25'd5535;
            NN[152]=25'd10342;
            NN[153]=25'd7411;
            NN[154]=25'd5944;
            NN[155]=25'd6659;
            NN[156]=25'd2071;
            NN[157]=25'd1360;
            NN[158]=25'd1503;
            NN[159]=25'd2747;
            NN[160]=25'd7743;
            NN[161]=25'd5903;
            NN[162]=25'd7036;
            NN[163]=25'd9426;
            NN[164]=25'd7293;
            NN[165]=-25'd717;
            NN[166]=-25'd584;
            NN[167]=-25'd66;
            NN[168]=25'd0;
            NN[169]=-25'd16;
            NN[170]=-25'd342;
            NN[171]=-25'd782;
            NN[172]=25'd2682;
            NN[173]=25'd16354;
            NN[174]=25'd18988;
            NN[175]=25'd9934;
            NN[176]=25'd23029;
            NN[177]=25'd22639;
            NN[178]=25'd8862;
            NN[179]=25'd16174;
            NN[180]=25'd9132;
            NN[181]=25'd5139;
            NN[182]=-25'd195;
            NN[183]=25'd2602;
            NN[184]=25'd6682;
            NN[185]=25'd6921;
            NN[186]=25'd4695;
            NN[187]=25'd4747;
            NN[188]=25'd3758;
            NN[189]=25'd10214;
            NN[190]=25'd18509;
            NN[191]=25'd10731;
            NN[192]=25'd3736;
            NN[193]=25'd796;
            NN[194]=-25'd105;
            NN[195]=25'd2;
            NN[196]=25'd0;
            NN[197]=-25'd7;
            NN[198]=-25'd459;
            NN[199]=25'd31;
            NN[200]=25'd4004;
            NN[201]=25'd2557;
            NN[202]=25'd5496;
            NN[203]=25'd11695;
            NN[204]=25'd16753;
            NN[205]=25'd16021;
            NN[206]=25'd8787;
            NN[207]=25'd8639;
            NN[208]=25'd6282;
            NN[209]=25'd1110;
            NN[210]=25'd3550;
            NN[211]=25'd6036;
            NN[212]=25'd5744;
            NN[213]=25'd7344;
            NN[214]=25'd738;
            NN[215]=25'd1282;
            NN[216]=25'd13879;
            NN[217]=25'd20775;
            NN[218]=25'd16609;
            NN[219]=25'd8750;
            NN[220]=25'd1832;
            NN[221]=25'd1256;
            NN[222]=25'd49;
            NN[223]=25'd0;
            NN[224]=25'd0;
            NN[225]=25'd0;
            NN[226]=-25'd395;
            NN[227]=25'd91;
            NN[228]=25'd4790;
            NN[229]=-25'd2765;
            NN[230]=-25'd7401;
            NN[231]=25'd345;
            NN[232]=25'd6255;
            NN[233]=25'd7879;
            NN[234]=25'd2065;
            NN[235]=25'd4874;
            NN[236]=25'd9866;
            NN[237]=25'd15082;
            NN[238]=25'd9244;
            NN[239]=25'd5896;
            NN[240]=25'd10142;
            NN[241]=25'd3937;
            NN[242]=25'd5511;
            NN[243]=25'd9299;
            NN[244]=25'd13965;
            NN[245]=25'd10770;
            NN[246]=25'd7817;
            NN[247]=25'd5555;
            NN[248]=25'd1818;
            NN[249]=25'd1281;
            NN[250]=25'd374;
            NN[251]=25'd0;
            NN[252]=25'd0;
            NN[253]=25'd0;
            NN[254]=-25'd81;
            NN[255]=25'd353;
            NN[256]=25'd2746;
            NN[257]=25'd1106;
            NN[258]=-25'd3935;
            NN[259]=-25'd5896;
            NN[260]=25'd2641;
            NN[261]=25'd8949;
            NN[262]=25'd14931;
            NN[263]=25'd12353;
            NN[264]=25'd13409;
            NN[265]=25'd6344;
            NN[266]=25'd7977;
            NN[267]=25'd3828;
            NN[268]=25'd7979;
            NN[269]=25'd614;
            NN[270]=-25'd2325;
            NN[271]=25'd4153;
            NN[272]=25'd7238;
            NN[273]=25'd2194;
            NN[274]=25'd2062;
            NN[275]=25'd2981;
            NN[276]=25'd1766;
            NN[277]=25'd900;
            NN[278]=25'd218;
            NN[279]=25'd0;
            NN[280]=25'd0;
            NN[281]=25'd0;
            NN[282]=-25'd23;
            NN[283]=25'd393;
            NN[284]=-25'd716;
            NN[285]=-25'd1845;
            NN[286]=-25'd1513;
            NN[287]=25'd990;
            NN[288]=25'd1639;
            NN[289]=25'd11193;
            NN[290]=25'd10658;
            NN[291]=25'd11525;
            NN[292]=25'd15049;
            NN[293]=25'd20161;
            NN[294]=25'd17015;
            NN[295]=25'd13085;
            NN[296]=25'd5134;
            NN[297]=25'd6581;
            NN[298]=25'd4225;
            NN[299]=25'd361;
            NN[300]=25'd142;
            NN[301]=-25'd36;
            NN[302]=25'd2133;
            NN[303]=25'd1919;
            NN[304]=25'd1350;
            NN[305]=-25'd200;
            NN[306]=-25'd6;
            NN[307]=25'd0;
            NN[308]=25'd0;
            NN[309]=25'd0;
            NN[310]=25'd0;
            NN[311]=25'd520;
            NN[312]=25'd287;
            NN[313]=-25'd1351;
            NN[314]=-25'd1582;
            NN[315]=-25'd847;
            NN[316]=25'd119;
            NN[317]=25'd4462;
            NN[318]=25'd6507;
            NN[319]=25'd10205;
            NN[320]=25'd11207;
            NN[321]=25'd11794;
            NN[322]=25'd7184;
            NN[323]=25'd9262;
            NN[324]=25'd7712;
            NN[325]=25'd6051;
            NN[326]=25'd1586;
            NN[327]=25'd900;
            NN[328]=25'd428;
            NN[329]=25'd1956;
            NN[330]=25'd2664;
            NN[331]=25'd1922;
            NN[332]=25'd1242;
            NN[333]=25'd0;
            NN[334]=25'd0;
            NN[335]=25'd0;
            NN[336]=25'd0;
            NN[337]=25'd0;
            NN[338]=25'd0;
            NN[339]=25'd0;
            NN[340]=-25'd230;
            NN[341]=-25'd466;
            NN[342]=-25'd691;
            NN[343]=-25'd1926;
            NN[344]=-25'd2404;
            NN[345]=-25'd1770;
            NN[346]=-25'd1127;
            NN[347]=25'd906;
            NN[348]=25'd1102;
            NN[349]=-25'd8;
            NN[350]=-25'd1982;
            NN[351]=25'd72;
            NN[352]=-25'd995;
            NN[353]=-25'd1439;
            NN[354]=-25'd2347;
            NN[355]=-25'd1305;
            NN[356]=25'd207;
            NN[357]=25'd333;
            NN[358]=25'd76;
            NN[359]=-25'd13;
            NN[360]=25'd0;
            NN[361]=25'd0;
            NN[362]=25'd0;
            NN[363]=25'd0;
            NN[364]=25'd0;
            NN[365]=25'd0;
            NN[366]=25'd0;
            NN[367]=25'd0;
            NN[368]=25'd0;
            NN[369]=25'd0;
            NN[370]=-25'd2;
            NN[371]=-25'd21;
            NN[372]=-25'd76;
            NN[373]=-25'd89;
            NN[374]=-25'd21;
            NN[375]=25'd41;
            NN[376]=-25'd54;
            NN[377]=-25'd251;
            NN[378]=-25'd493;
            NN[379]=-25'd402;
            NN[380]=-25'd424;
            NN[381]=-25'd427;
            NN[382]=-25'd336;
            NN[383]=-25'd270;
            NN[384]=-25'd284;
            NN[385]=-25'd103;
            NN[386]=-25'd74;
            NN[387]=-25'd16;
            NN[388]=25'd0;
            NN[389]=25'd0;
            NN[390]=25'd0;
            NN[391]=25'd0;
        end
        12:begin
            NN[0]=25'd0;
            NN[1]=25'd0;
            NN[2]=25'd0;
            NN[3]=25'd0;
            NN[4]=25'd0;
            NN[5]=25'd0;
            NN[6]=25'd0;
            NN[7]=25'd0;
            NN[8]=25'd0;
            NN[9]=25'd0;
            NN[10]=25'd0;
            NN[11]=25'd0;
            NN[12]=25'd217;
            NN[13]=25'd475;
            NN[14]=25'd0;
            NN[15]=25'd0;
            NN[16]=25'd0;
            NN[17]=25'd0;
            NN[18]=25'd0;
            NN[19]=25'd0;
            NN[20]=25'd0;
            NN[21]=25'd0;
            NN[22]=25'd0;
            NN[23]=25'd0;
            NN[24]=25'd0;
            NN[25]=25'd0;
            NN[26]=25'd0;
            NN[27]=25'd0;
            NN[28]=25'd0;
            NN[29]=25'd0;
            NN[30]=25'd0;
            NN[31]=25'd0;
            NN[32]=25'd2;
            NN[33]=25'd9;
            NN[34]=25'd616;
            NN[35]=25'd1461;
            NN[36]=25'd1772;
            NN[37]=25'd1495;
            NN[38]=25'd3124;
            NN[39]=25'd3098;
            NN[40]=25'd4978;
            NN[41]=25'd3132;
            NN[42]=25'd1202;
            NN[43]=25'd1080;
            NN[44]=25'd1242;
            NN[45]=25'd1238;
            NN[46]=25'd1257;
            NN[47]=25'd948;
            NN[48]=25'd673;
            NN[49]=25'd776;
            NN[50]=25'd687;
            NN[51]=25'd201;
            NN[52]=25'd0;
            NN[53]=25'd0;
            NN[54]=25'd0;
            NN[55]=25'd0;
            NN[56]=25'd0;
            NN[57]=25'd0;
            NN[58]=25'd0;
            NN[59]=25'd4;
            NN[60]=25'd35;
            NN[61]=25'd36;
            NN[62]=25'd912;
            NN[63]=25'd3318;
            NN[64]=25'd5231;
            NN[65]=25'd7204;
            NN[66]=25'd12483;
            NN[67]=25'd13609;
            NN[68]=25'd17252;
            NN[69]=25'd14777;
            NN[70]=25'd12032;
            NN[71]=25'd10165;
            NN[72]=25'd12011;
            NN[73]=25'd10436;
            NN[74]=25'd9687;
            NN[75]=25'd9191;
            NN[76]=25'd7223;
            NN[77]=25'd6903;
            NN[78]=25'd5492;
            NN[79]=25'd2269;
            NN[80]=-25'd52;
            NN[81]=-25'd321;
            NN[82]=25'd0;
            NN[83]=25'd0;
            NN[84]=25'd0;
            NN[85]=25'd0;
            NN[86]=-25'd4;
            NN[87]=25'd57;
            NN[88]=25'd116;
            NN[89]=25'd331;
            NN[90]=25'd2125;
            NN[91]=25'd4175;
            NN[92]=25'd6842;
            NN[93]=25'd9628;
            NN[94]=25'd12381;
            NN[95]=25'd14605;
            NN[96]=25'd12591;
            NN[97]=25'd14237;
            NN[98]=25'd16446;
            NN[99]=25'd16607;
            NN[100]=25'd15505;
            NN[101]=25'd14530;
            NN[102]=25'd18766;
            NN[103]=25'd21536;
            NN[104]=25'd17407;
            NN[105]=25'd16812;
            NN[106]=25'd13677;
            NN[107]=25'd9532;
            NN[108]=25'd5066;
            NN[109]=-25'd169;
            NN[110]=25'd355;
            NN[111]=25'd0;
            NN[112]=25'd0;
            NN[113]=25'd0;
            NN[114]=-25'd18;
            NN[115]=-25'd63;
            NN[116]=25'd117;
            NN[117]=-25'd314;
            NN[118]=-25'd389;
            NN[119]=25'd1958;
            NN[120]=25'd5878;
            NN[121]=25'd4507;
            NN[122]=25'd5093;
            NN[123]=-25'd620;
            NN[124]=-25'd2160;
            NN[125]=-25'd562;
            NN[126]=-25'd999;
            NN[127]=-25'd1774;
            NN[128]=25'd3949;
            NN[129]=25'd12145;
            NN[130]=25'd16123;
            NN[131]=25'd21722;
            NN[132]=25'd21769;
            NN[133]=25'd20566;
            NN[134]=25'd18185;
            NN[135]=25'd11726;
            NN[136]=25'd3789;
            NN[137]=25'd654;
            NN[138]=25'd1;
            NN[139]=25'd237;
            NN[140]=25'd0;
            NN[141]=25'd0;
            NN[142]=25'd0;
            NN[143]=-25'd669;
            NN[144]=-25'd179;
            NN[145]=-25'd3589;
            NN[146]=-25'd2886;
            NN[147]=-25'd1560;
            NN[148]=25'd2545;
            NN[149]=25'd770;
            NN[150]=-25'd1525;
            NN[151]=-25'd13138;
            NN[152]=-25'd11452;
            NN[153]=-25'd14602;
            NN[154]=-25'd8584;
            NN[155]=-25'd10238;
            NN[156]=-25'd6456;
            NN[157]=25'd1647;
            NN[158]=25'd9883;
            NN[159]=25'd14608;
            NN[160]=25'd13173;
            NN[161]=25'd9930;
            NN[162]=25'd7352;
            NN[163]=25'd7699;
            NN[164]=25'd3015;
            NN[165]=-25'd504;
            NN[166]=25'd465;
            NN[167]=25'd354;
            NN[168]=25'd0;
            NN[169]=25'd0;
            NN[170]=-25'd19;
            NN[171]=-25'd1061;
            NN[172]=-25'd973;
            NN[173]=-25'd3865;
            NN[174]=-25'd6149;
            NN[175]=-25'd1803;
            NN[176]=-25'd1080;
            NN[177]=-25'd4859;
            NN[178]=-25'd13396;
            NN[179]=-25'd14986;
            NN[180]=-25'd11624;
            NN[181]=-25'd14781;
            NN[182]=-25'd16188;
            NN[183]=-25'd12987;
            NN[184]=-25'd14091;
            NN[185]=-25'd10581;
            NN[186]=-25'd10519;
            NN[187]=-25'd6058;
            NN[188]=-25'd4585;
            NN[189]=-25'd3926;
            NN[190]=-25'd4711;
            NN[191]=-25'd5087;
            NN[192]=-25'd3683;
            NN[193]=-25'd2152;
            NN[194]=-25'd1127;
            NN[195]=-25'd86;
            NN[196]=25'd0;
            NN[197]=25'd0;
            NN[198]=-25'd143;
            NN[199]=-25'd1441;
            NN[200]=-25'd1613;
            NN[201]=-25'd4327;
            NN[202]=-25'd7425;
            NN[203]=-25'd1518;
            NN[204]=-25'd2125;
            NN[205]=-25'd8365;
            NN[206]=-25'd14468;
            NN[207]=-25'd14004;
            NN[208]=-25'd14104;
            NN[209]=-25'd18131;
            NN[210]=-25'd17367;
            NN[211]=-25'd15297;
            NN[212]=-25'd21289;
            NN[213]=-25'd22649;
            NN[214]=-25'd25643;
            NN[215]=-25'd24514;
            NN[216]=-25'd21307;
            NN[217]=-25'd18464;
            NN[218]=-25'd19106;
            NN[219]=-25'd15271;
            NN[220]=-25'd6720;
            NN[221]=-25'd4273;
            NN[222]=-25'd1173;
            NN[223]=-25'd211;
            NN[224]=25'd0;
            NN[225]=-25'd12;
            NN[226]=-25'd206;
            NN[227]=-25'd1665;
            NN[228]=-25'd2203;
            NN[229]=-25'd6291;
            NN[230]=-25'd8414;
            NN[231]=-25'd5007;
            NN[232]=-25'd5559;
            NN[233]=-25'd10311;
            NN[234]=-25'd13575;
            NN[235]=-25'd15406;
            NN[236]=-25'd16712;
            NN[237]=-25'd19469;
            NN[238]=-25'd21479;
            NN[239]=-25'd24636;
            NN[240]=-25'd31825;
            NN[241]=-25'd37115;
            NN[242]=-25'd43610;
            NN[243]=-25'd39576;
            NN[244]=-25'd30885;
            NN[245]=-25'd26647;
            NN[246]=-25'd26398;
            NN[247]=-25'd19937;
            NN[248]=-25'd12374;
            NN[249]=-25'd5966;
            NN[250]=-25'd2516;
            NN[251]=-25'd133;
            NN[252]=25'd0;
            NN[253]=-25'd1;
            NN[254]=-25'd246;
            NN[255]=-25'd2128;
            NN[256]=-25'd2866;
            NN[257]=-25'd8177;
            NN[258]=-25'd8106;
            NN[259]=-25'd1850;
            NN[260]=-25'd2325;
            NN[261]=-25'd10130;
            NN[262]=-25'd12672;
            NN[263]=-25'd11612;
            NN[264]=-25'd13862;
            NN[265]=-25'd19014;
            NN[266]=-25'd13793;
            NN[267]=-25'd27630;
            NN[268]=-25'd41284;
            NN[269]=-25'd48464;
            NN[270]=-25'd46884;
            NN[271]=-25'd40392;
            NN[272]=-25'd30949;
            NN[273]=-25'd25452;
            NN[274]=-25'd26527;
            NN[275]=-25'd16591;
            NN[276]=-25'd12550;
            NN[277]=-25'd9303;
            NN[278]=-25'd3385;
            NN[279]=-25'd191;
            NN[280]=25'd0;
            NN[281]=-25'd1;
            NN[282]=-25'd550;
            NN[283]=-25'd2122;
            NN[284]=-25'd3444;
            NN[285]=-25'd6965;
            NN[286]=-25'd4422;
            NN[287]=25'd3856;
            NN[288]=25'd2378;
            NN[289]=-25'd5717;
            NN[290]=-25'd4247;
            NN[291]=-25'd4602;
            NN[292]=-25'd10202;
            NN[293]=-25'd6560;
            NN[294]=-25'd15555;
            NN[295]=-25'd33410;
            NN[296]=-25'd39653;
            NN[297]=-25'd39920;
            NN[298]=-25'd35910;
            NN[299]=-25'd30775;
            NN[300]=-25'd23305;
            NN[301]=-25'd18281;
            NN[302]=-25'd15242;
            NN[303]=-25'd7750;
            NN[304]=-25'd9826;
            NN[305]=-25'd10629;
            NN[306]=-25'd3117;
            NN[307]=-25'd475;
            NN[308]=25'd0;
            NN[309]=-25'd21;
            NN[310]=-25'd76;
            NN[311]=-25'd1878;
            NN[312]=-25'd2366;
            NN[313]=-25'd710;
            NN[314]=25'd1705;
            NN[315]=25'd9834;
            NN[316]=25'd5189;
            NN[317]=25'd6422;
            NN[318]=25'd4576;
            NN[319]=25'd1050;
            NN[320]=25'd5991;
            NN[321]=25'd5392;
            NN[322]=-25'd17863;
            NN[323]=-25'd36769;
            NN[324]=-25'd26963;
            NN[325]=-25'd23070;
            NN[326]=-25'd18845;
            NN[327]=-25'd15761;
            NN[328]=-25'd8719;
            NN[329]=-25'd75;
            NN[330]=25'd5422;
            NN[331]=25'd11004;
            NN[332]=-25'd889;
            NN[333]=-25'd8163;
            NN[334]=-25'd3658;
            NN[335]=-25'd297;
            NN[336]=25'd0;
            NN[337]=-25'd31;
            NN[338]=-25'd68;
            NN[339]=-25'd1481;
            NN[340]=-25'd2827;
            NN[341]=25'd1631;
            NN[342]=25'd10888;
            NN[343]=25'd13361;
            NN[344]=25'd9683;
            NN[345]=25'd12160;
            NN[346]=25'd6375;
            NN[347]=25'd15222;
            NN[348]=25'd15227;
            NN[349]=25'd6377;
            NN[350]=-25'd20046;
            NN[351]=-25'd21271;
            NN[352]=-25'd7695;
            NN[353]=-25'd8517;
            NN[354]=-25'd9319;
            NN[355]=-25'd11919;
            NN[356]=-25'd2192;
            NN[357]=25'd11445;
            NN[358]=25'd21419;
            NN[359]=25'd28380;
            NN[360]=25'd11859;
            NN[361]=-25'd4261;
            NN[362]=-25'd3276;
            NN[363]=-25'd162;
            NN[364]=25'd0;
            NN[365]=-25'd33;
            NN[366]=-25'd25;
            NN[367]=-25'd1232;
            NN[368]=-25'd3651;
            NN[369]=25'd4936;
            NN[370]=25'd17306;
            NN[371]=25'd10267;
            NN[372]=25'd9774;
            NN[373]=25'd11297;
            NN[374]=25'd15473;
            NN[375]=25'd17794;
            NN[376]=25'd11769;
            NN[377]=-25'd2565;
            NN[378]=-25'd13354;
            NN[379]=25'd2363;
            NN[380]=25'd5325;
            NN[381]=-25'd6457;
            NN[382]=-25'd11917;
            NN[383]=-25'd4336;
            NN[384]=25'd935;
            NN[385]=25'd17696;
            NN[386]=25'd29024;
            NN[387]=25'd35556;
            NN[388]=25'd18509;
            NN[389]=-25'd4321;
            NN[390]=-25'd3954;
            NN[391]=-25'd530;
        end
        13:begin
            NN[0]=-25'd8;
            NN[1]=-25'd2;
            NN[2]=-25'd6;
            NN[3]=-25'd936;
            NN[4]=-25'd7114;
            NN[5]=25'd3392;
            NN[6]=25'd13891;
            NN[7]=25'd10509;
            NN[8]=25'd12089;
            NN[9]=25'd15961;
            NN[10]=25'd21913;
            NN[11]=25'd27943;
            NN[12]=25'd11085;
            NN[13]=-25'd8182;
            NN[14]=-25'd2449;
            NN[15]=25'd6984;
            NN[16]=25'd6960;
            NN[17]=-25'd12984;
            NN[18]=-25'd11865;
            NN[19]=-25'd4164;
            NN[20]=25'd1149;
            NN[21]=25'd15031;
            NN[22]=25'd27292;
            NN[23]=25'd29942;
            NN[24]=25'd14383;
            NN[25]=-25'd3367;
            NN[26]=-25'd4146;
            NN[27]=-25'd84;
            NN[28]=-25'd2;
            NN[29]=-25'd4;
            NN[30]=-25'd22;
            NN[31]=-25'd2465;
            NN[32]=-25'd11189;
            NN[33]=-25'd889;
            NN[34]=25'd11429;
            NN[35]=25'd15439;
            NN[36]=25'd15613;
            NN[37]=25'd17322;
            NN[38]=25'd31466;
            NN[39]=25'd32763;
            NN[40]=25'd10783;
            NN[41]=25'd2854;
            NN[42]=25'd13671;
            NN[43]=25'd10231;
            NN[44]=25'd822;
            NN[45]=-25'd9787;
            NN[46]=-25'd8769;
            NN[47]=25'd312;
            NN[48]=25'd8556;
            NN[49]=25'd16357;
            NN[50]=25'd15344;
            NN[51]=25'd17852;
            NN[52]=25'd8577;
            NN[53]=-25'd3142;
            NN[54]=-25'd4972;
            NN[55]=-25'd435;
            NN[56]=25'd0;
            NN[57]=-25'd2;
            NN[58]=-25'd89;
            NN[59]=-25'd4036;
            NN[60]=-25'd13707;
            NN[61]=-25'd4314;
            NN[62]=25'd10227;
            NN[63]=25'd19205;
            NN[64]=25'd20285;
            NN[65]=25'd24780;
            NN[66]=25'd38049;
            NN[67]=25'd39076;
            NN[68]=25'd7631;
            NN[69]=25'd6129;
            NN[70]=25'd15005;
            NN[71]=25'd9118;
            NN[72]=-25'd6530;
            NN[73]=-25'd11822;
            NN[74]=25'd707;
            NN[75]=25'd7985;
            NN[76]=25'd6709;
            NN[77]=25'd5830;
            NN[78]=25'd4494;
            NN[79]=25'd5962;
            NN[80]=25'd2402;
            NN[81]=-25'd5706;
            NN[82]=-25'd4534;
            NN[83]=-25'd676;
            NN[84]=25'd0;
            NN[85]=-25'd1;
            NN[86]=-25'd187;
            NN[87]=-25'd4713;
            NN[88]=-25'd16943;
            NN[89]=-25'd10131;
            NN[90]=25'd2096;
            NN[91]=25'd16328;
            NN[92]=25'd21315;
            NN[93]=25'd23538;
            NN[94]=25'd41241;
            NN[95]=25'd39916;
            NN[96]=25'd15857;
            NN[97]=25'd8460;
            NN[98]=25'd10625;
            NN[99]=25'd1754;
            NN[100]=-25'd8243;
            NN[101]=25'd2002;
            NN[102]=25'd12907;
            NN[103]=25'd13569;
            NN[104]=25'd7401;
            NN[105]=25'd5372;
            NN[106]=25'd3190;
            NN[107]=25'd718;
            NN[108]=-25'd4039;
            NN[109]=-25'd5637;
            NN[110]=-25'd3010;
            NN[111]=-25'd362;
            NN[112]=-25'd3;
            NN[113]=25'd0;
            NN[114]=-25'd135;
            NN[115]=-25'd4795;
            NN[116]=-25'd16328;
            NN[117]=-25'd18740;
            NN[118]=-25'd6015;
            NN[119]=25'd12442;
            NN[120]=25'd18057;
            NN[121]=25'd20719;
            NN[122]=25'd31641;
            NN[123]=25'd35790;
            NN[124]=25'd33079;
            NN[125]=25'd16325;
            NN[126]=25'd6828;
            NN[127]=25'd6376;
            NN[128]=25'd11418;
            NN[129]=25'd17284;
            NN[130]=25'd18606;
            NN[131]=25'd8494;
            NN[132]=25'd6554;
            NN[133]=25'd5838;
            NN[134]=25'd2605;
            NN[135]=-25'd1342;
            NN[136]=-25'd6048;
            NN[137]=-25'd2841;
            NN[138]=-25'd783;
            NN[139]=-25'd448;
            NN[140]=25'd0;
            NN[141]=-25'd20;
            NN[142]=-25'd160;
            NN[143]=-25'd4693;
            NN[144]=-25'd13798;
            NN[145]=-25'd19530;
            NN[146]=-25'd12103;
            NN[147]=25'd5183;
            NN[148]=25'd10765;
            NN[149]=25'd17902;
            NN[150]=25'd32280;
            NN[151]=25'd44533;
            NN[152]=25'd40549;
            NN[153]=25'd21731;
            NN[154]=25'd18416;
            NN[155]=25'd18632;
            NN[156]=25'd21802;
            NN[157]=25'd18053;
            NN[158]=25'd13576;
            NN[159]=25'd12814;
            NN[160]=25'd9830;
            NN[161]=25'd5687;
            NN[162]=25'd1069;
            NN[163]=-25'd4948;
            NN[164]=-25'd5935;
            NN[165]=-25'd4419;
            NN[166]=-25'd1535;
            NN[167]=-25'd308;
            NN[168]=25'd0;
            NN[169]=-25'd44;
            NN[170]=-25'd158;
            NN[171]=-25'd3344;
            NN[172]=-25'd11441;
            NN[173]=-25'd19854;
            NN[174]=-25'd18932;
            NN[175]=-25'd3979;
            NN[176]=25'd343;
            NN[177]=25'd14746;
            NN[178]=25'd30253;
            NN[179]=25'd34279;
            NN[180]=25'd42096;
            NN[181]=25'd34063;
            NN[182]=25'd37857;
            NN[183]=25'd29033;
            NN[184]=25'd21627;
            NN[185]=25'd13832;
            NN[186]=25'd17411;
            NN[187]=25'd10089;
            NN[188]=25'd7969;
            NN[189]=-25'd1014;
            NN[190]=-25'd7845;
            NN[191]=-25'd5101;
            NN[192]=-25'd4411;
            NN[193]=-25'd1858;
            NN[194]=-25'd412;
            NN[195]=25'd0;
            NN[196]=25'd0;
            NN[197]=25'd0;
            NN[198]=-25'd72;
            NN[199]=-25'd1369;
            NN[200]=-25'd7600;
            NN[201]=-25'd15419;
            NN[202]=-25'd22373;
            NN[203]=-25'd14726;
            NN[204]=-25'd3307;
            NN[205]=25'd5182;
            NN[206]=25'd17219;
            NN[207]=25'd27745;
            NN[208]=25'd40814;
            NN[209]=25'd43812;
            NN[210]=25'd39636;
            NN[211]=25'd26553;
            NN[212]=25'd18659;
            NN[213]=25'd18106;
            NN[214]=25'd13605;
            NN[215]=25'd5045;
            NN[216]=-25'd1383;
            NN[217]=-25'd6109;
            NN[218]=-25'd4740;
            NN[219]=-25'd3151;
            NN[220]=-25'd1672;
            NN[221]=-25'd729;
            NN[222]=-25'd103;
            NN[223]=25'd0;
            NN[224]=25'd0;
            NN[225]=25'd0;
            NN[226]=-25'd18;
            NN[227]=-25'd294;
            NN[228]=-25'd3325;
            NN[229]=-25'd8646;
            NN[230]=-25'd16449;
            NN[231]=-25'd20518;
            NN[232]=-25'd19890;
            NN[233]=-25'd14032;
            NN[234]=-25'd7367;
            NN[235]=-25'd1022;
            NN[236]=25'd9290;
            NN[237]=25'd8908;
            NN[238]=25'd4424;
            NN[239]=25'd5299;
            NN[240]=25'd2540;
            NN[241]=-25'd1104;
            NN[242]=-25'd6712;
            NN[243]=-25'd7446;
            NN[244]=-25'd5313;
            NN[245]=-25'd4318;
            NN[246]=-25'd5535;
            NN[247]=-25'd3342;
            NN[248]=-25'd1118;
            NN[249]=-25'd314;
            NN[250]=-25'd8;
            NN[251]=25'd0;
            NN[252]=25'd0;
            NN[253]=25'd0;
            NN[254]=-25'd3;
            NN[255]=-25'd103;
            NN[256]=-25'd860;
            NN[257]=-25'd2750;
            NN[258]=-25'd6399;
            NN[259]=-25'd13034;
            NN[260]=-25'd19329;
            NN[261]=-25'd23496;
            NN[262]=-25'd28213;
            NN[263]=-25'd27864;
            NN[264]=-25'd21733;
            NN[265]=-25'd16656;
            NN[266]=-25'd13709;
            NN[267]=-25'd12009;
            NN[268]=-25'd12988;
            NN[269]=-25'd12934;
            NN[270]=-25'd8970;
            NN[271]=-25'd6773;
            NN[272]=-25'd6061;
            NN[273]=-25'd5007;
            NN[274]=-25'd2982;
            NN[275]=-25'd1548;
            NN[276]=-25'd646;
            NN[277]=-25'd143;
            NN[278]=-25'd7;
            NN[279]=25'd0;
            NN[280]=25'd0;
            NN[281]=25'd0;
            NN[282]=25'd0;
            NN[283]=-25'd4;
            NN[284]=-25'd148;
            NN[285]=-25'd698;
            NN[286]=-25'd1528;
            NN[287]=-25'd3680;
            NN[288]=-25'd7124;
            NN[289]=-25'd10754;
            NN[290]=-25'd13728;
            NN[291]=-25'd17287;
            NN[292]=-25'd17963;
            NN[293]=-25'd18890;
            NN[294]=-25'd17788;
            NN[295]=-25'd16301;
            NN[296]=-25'd13001;
            NN[297]=-25'd9738;
            NN[298]=-25'd7086;
            NN[299]=-25'd5467;
            NN[300]=-25'd3497;
            NN[301]=-25'd2616;
            NN[302]=-25'd1451;
            NN[303]=-25'd571;
            NN[304]=-25'd118;
            NN[305]=-25'd16;
            NN[306]=-25'd1;
            NN[307]=25'd0;
            NN[308]=25'd0;
            NN[309]=25'd0;
            NN[310]=25'd0;
            NN[311]=-25'd1;
            NN[312]=-25'd47;
            NN[313]=-25'd156;
            NN[314]=-25'd471;
            NN[315]=-25'd1020;
            NN[316]=-25'd2286;
            NN[317]=-25'd3034;
            NN[318]=-25'd3186;
            NN[319]=-25'd3774;
            NN[320]=-25'd4446;
            NN[321]=-25'd5555;
            NN[322]=-25'd5443;
            NN[323]=-25'd5118;
            NN[324]=-25'd4236;
            NN[325]=-25'd3085;
            NN[326]=-25'd2311;
            NN[327]=-25'd1709;
            NN[328]=-25'd956;
            NN[329]=-25'd541;
            NN[330]=-25'd259;
            NN[331]=-25'd132;
            NN[332]=-25'd25;
            NN[333]=-25'd1;
            NN[334]=-25'd1;
            NN[335]=25'd0;
            NN[336]=25'd0;
            NN[337]=25'd0;
            NN[338]=25'd0;
            NN[339]=25'd0;
            NN[340]=-25'd8;
            NN[341]=-25'd17;
            NN[342]=-25'd51;
            NN[343]=-25'd142;
            NN[344]=-25'd239;
            NN[345]=-25'd348;
            NN[346]=-25'd568;
            NN[347]=-25'd868;
            NN[348]=-25'd961;
            NN[349]=-25'd1201;
            NN[350]=-25'd1009;
            NN[351]=-25'd991;
            NN[352]=-25'd1035;
            NN[353]=-25'd775;
            NN[354]=-25'd563;
            NN[355]=-25'd327;
            NN[356]=-25'd145;
            NN[357]=-25'd78;
            NN[358]=-25'd31;
            NN[359]=-25'd4;
            NN[360]=25'd0;
            NN[361]=25'd0;
            NN[362]=25'd0;
            NN[363]=25'd0;
            NN[364]=25'd0;
            NN[365]=25'd0;
            NN[366]=25'd0;
            NN[367]=25'd0;
            NN[368]=25'd0;
            NN[369]=25'd0;
            NN[370]=25'd0;
            NN[371]=-25'd4;
            NN[372]=-25'd9;
            NN[373]=-25'd14;
            NN[374]=-25'd32;
            NN[375]=-25'd65;
            NN[376]=-25'd80;
            NN[377]=-25'd92;
            NN[378]=-25'd102;
            NN[379]=-25'd81;
            NN[380]=-25'd98;
            NN[381]=-25'd80;
            NN[382]=-25'd29;
            NN[383]=-25'd7;
            NN[384]=-25'd7;
            NN[385]=-25'd5;
            NN[386]=-25'd10;
            NN[387]=-25'd2;
            NN[388]=25'd0;
            NN[389]=25'd0;
            NN[390]=25'd0;
            NN[391]=25'd0;
        end
        14:begin
            NN[0]=25'd0;
            NN[1]=25'd0;
            NN[2]=25'd0;
            NN[3]=25'd0;
            NN[4]=25'd0;
            NN[5]=25'd0;
            NN[6]=25'd0;
            NN[7]=25'd0;
            NN[8]=25'd0;
            NN[9]=25'd0;
            NN[10]=25'd0;
            NN[11]=25'd0;
            NN[12]=25'd0;
            NN[13]=25'd0;
            NN[14]=25'd0;
            NN[15]=25'd0;
            NN[16]=25'd0;
            NN[17]=25'd0;
            NN[18]=25'd0;
            NN[19]=25'd0;
            NN[20]=25'd0;
            NN[21]=25'd0;
            NN[22]=25'd0;
            NN[23]=25'd0;
            NN[24]=25'd0;
            NN[25]=25'd0;
            NN[26]=25'd0;
            NN[27]=25'd0;
            NN[28]=25'd0;
            NN[29]=25'd0;
            NN[30]=25'd0;
            NN[31]=25'd0;
            NN[32]=25'd0;
            NN[33]=25'd0;
            NN[34]=-25'd1;
            NN[35]=-25'd8;
            NN[36]=-25'd51;
            NN[37]=-25'd95;
            NN[38]=-25'd177;
            NN[39]=-25'd248;
            NN[40]=-25'd397;
            NN[41]=-25'd140;
            NN[42]=-25'd18;
            NN[43]=-25'd63;
            NN[44]=-25'd172;
            NN[45]=-25'd45;
            NN[46]=-25'd9;
            NN[47]=-25'd20;
            NN[48]=-25'd11;
            NN[49]=25'd0;
            NN[50]=25'd0;
            NN[51]=25'd0;
            NN[52]=25'd0;
            NN[53]=25'd0;
            NN[54]=25'd0;
            NN[55]=25'd0;
            NN[56]=25'd0;
            NN[57]=25'd0;
            NN[58]=25'd0;
            NN[59]=-25'd2;
            NN[60]=-25'd1;
            NN[61]=25'd0;
            NN[62]=-25'd13;
            NN[63]=-25'd68;
            NN[64]=-25'd212;
            NN[65]=-25'd450;
            NN[66]=-25'd742;
            NN[67]=-25'd1120;
            NN[68]=-25'd958;
            NN[69]=-25'd577;
            NN[70]=-25'd630;
            NN[71]=-25'd801;
            NN[72]=-25'd660;
            NN[73]=-25'd458;
            NN[74]=-25'd292;
            NN[75]=-25'd169;
            NN[76]=-25'd100;
            NN[77]=-25'd110;
            NN[78]=-25'd84;
            NN[79]=-25'd6;
            NN[80]=25'd0;
            NN[81]=25'd0;
            NN[82]=25'd0;
            NN[83]=25'd0;
            NN[84]=25'd0;
            NN[85]=25'd0;
            NN[86]=25'd0;
            NN[87]=-25'd8;
            NN[88]=-25'd29;
            NN[89]=-25'd32;
            NN[90]=-25'd87;
            NN[91]=-25'd403;
            NN[92]=-25'd1223;
            NN[93]=-25'd1872;
            NN[94]=-25'd3073;
            NN[95]=-25'd3872;
            NN[96]=-25'd3210;
            NN[97]=-25'd3127;
            NN[98]=-25'd3276;
            NN[99]=-25'd3607;
            NN[100]=-25'd3166;
            NN[101]=-25'd2489;
            NN[102]=-25'd2170;
            NN[103]=-25'd1323;
            NN[104]=-25'd1024;
            NN[105]=-25'd628;
            NN[106]=-25'd276;
            NN[107]=-25'd124;
            NN[108]=-25'd44;
            NN[109]=-25'd1;
            NN[110]=25'd0;
            NN[111]=25'd0;
            NN[112]=25'd0;
            NN[113]=25'd0;
            NN[114]=25'd0;
            NN[115]=25'd26;
            NN[116]=-25'd76;
            NN[117]=-25'd581;
            NN[118]=-25'd751;
            NN[119]=-25'd1821;
            NN[120]=-25'd3287;
            NN[121]=-25'd5687;
            NN[122]=-25'd8426;
            NN[123]=-25'd10325;
            NN[124]=-25'd12075;
            NN[125]=-25'd14014;
            NN[126]=-25'd15824;
            NN[127]=-25'd15993;
            NN[128]=-25'd14739;
            NN[129]=-25'd12186;
            NN[130]=-25'd9640;
            NN[131]=-25'd6878;
            NN[132]=-25'd5347;
            NN[133]=-25'd3055;
            NN[134]=-25'd2080;
            NN[135]=-25'd971;
            NN[136]=-25'd382;
            NN[137]=-25'd101;
            NN[138]=-25'd29;
            NN[139]=-25'd1;
            NN[140]=25'd0;
            NN[141]=25'd0;
            NN[142]=25'd0;
            NN[143]=-25'd5;
            NN[144]=-25'd107;
            NN[145]=25'd1107;
            NN[146]=25'd1202;
            NN[147]=25'd65;
            NN[148]=-25'd816;
            NN[149]=-25'd5103;
            NN[150]=-25'd10811;
            NN[151]=-25'd16116;
            NN[152]=-25'd19612;
            NN[153]=-25'd26098;
            NN[154]=-25'd31399;
            NN[155]=-25'd33016;
            NN[156]=-25'd30356;
            NN[157]=-25'd28927;
            NN[158]=-25'd26629;
            NN[159]=-25'd23084;
            NN[160]=-25'd18701;
            NN[161]=-25'd11852;
            NN[162]=-25'd7674;
            NN[163]=-25'd4504;
            NN[164]=-25'd1850;
            NN[165]=-25'd668;
            NN[166]=-25'd250;
            NN[167]=-25'd11;
            NN[168]=25'd0;
            NN[169]=25'd0;
            NN[170]=25'd292;
            NN[171]=25'd1528;
            NN[172]=25'd1294;
            NN[173]=25'd3824;
            NN[174]=25'd7697;
            NN[175]=25'd8192;
            NN[176]=25'd10919;
            NN[177]=25'd7782;
            NN[178]=25'd9563;
            NN[179]=25'd7923;
            NN[180]=-25'd2390;
            NN[181]=-25'd12745;
            NN[182]=-25'd17092;
            NN[183]=-25'd12484;
            NN[184]=-25'd10332;
            NN[185]=-25'd10469;
            NN[186]=-25'd13181;
            NN[187]=-25'd12575;
            NN[188]=-25'd11295;
            NN[189]=-25'd6958;
            NN[190]=-25'd9285;
            NN[191]=-25'd8323;
            NN[192]=-25'd4932;
            NN[193]=-25'd2420;
            NN[194]=-25'd832;
            NN[195]=-25'd101;
            NN[196]=25'd0;
            NN[197]=25'd121;
            NN[198]=25'd1571;
            NN[199]=25'd4862;
            NN[200]=25'd4383;
            NN[201]=25'd8871;
            NN[202]=25'd15399;
            NN[203]=25'd17988;
            NN[204]=25'd19271;
            NN[205]=25'd20347;
            NN[206]=25'd24539;
            NN[207]=25'd23283;
            NN[208]=25'd18832;
            NN[209]=25'd11350;
            NN[210]=25'd929;
            NN[211]=25'd3201;
            NN[212]=25'd11682;
            NN[213]=25'd15610;
            NN[214]=25'd14098;
            NN[215]=25'd9636;
            NN[216]=25'd6803;
            NN[217]=25'd2212;
            NN[218]=25'd1415;
            NN[219]=-25'd2894;
            NN[220]=-25'd5437;
            NN[221]=-25'd3908;
            NN[222]=-25'd815;
            NN[223]=-25'd85;
            NN[224]=-25'd65;
            NN[225]=25'd1171;
            NN[226]=25'd3957;
            NN[227]=25'd9841;
            NN[228]=25'd12864;
            NN[229]=25'd15924;
            NN[230]=25'd16198;
            NN[231]=25'd22854;
            NN[232]=25'd16158;
            NN[233]=25'd12497;
            NN[234]=25'd14556;
            NN[235]=25'd23684;
            NN[236]=25'd24729;
            NN[237]=25'd13623;
            NN[238]=25'd17967;
            NN[239]=25'd23317;
            NN[240]=25'd26133;
            NN[241]=25'd24289;
            NN[242]=25'd25903;
            NN[243]=25'd16570;
            NN[244]=25'd12882;
            NN[245]=25'd4576;
            NN[246]=25'd5910;
            NN[247]=-25'd589;
            NN[248]=-25'd7074;
            NN[249]=-25'd4710;
            NN[250]=-25'd1289;
            NN[251]=-25'd234;
            NN[252]=25'd80;
            NN[253]=25'd1565;
            NN[254]=25'd4750;
            NN[255]=25'd13191;
            NN[256]=25'd18634;
            NN[257]=25'd15433;
            NN[258]=25'd10549;
            NN[259]=25'd8183;
            NN[260]=25'd4666;
            NN[261]=25'd5158;
            NN[262]=25'd4178;
            NN[263]=25'd11103;
            NN[264]=25'd15002;
            NN[265]=25'd14961;
            NN[266]=25'd25145;
            NN[267]=25'd33022;
            NN[268]=25'd36887;
            NN[269]=25'd35578;
            NN[270]=25'd25768;
            NN[271]=25'd24683;
            NN[272]=25'd14538;
            NN[273]=25'd14450;
            NN[274]=25'd7752;
            NN[275]=-25'd4950;
            NN[276]=-25'd7294;
            NN[277]=-25'd3546;
            NN[278]=-25'd655;
            NN[279]=25'd678;
            NN[280]=25'd102;
            NN[281]=25'd1556;
            NN[282]=25'd5499;
            NN[283]=25'd12256;
            NN[284]=25'd18160;
            NN[285]=25'd15623;
            NN[286]=25'd5624;
            NN[287]=25'd3047;
            NN[288]=-25'd4157;
            NN[289]=25'd3391;
            NN[290]=25'd5656;
            NN[291]=25'd1042;
            NN[292]=25'd482;
            NN[293]=25'd15843;
            NN[294]=25'd26748;
            NN[295]=25'd40481;
            NN[296]=25'd49149;
            NN[297]=25'd38083;
            NN[298]=25'd27945;
            NN[299]=25'd24993;
            NN[300]=25'd22249;
            NN[301]=25'd20606;
            NN[302]=25'd8980;
            NN[303]=-25'd8224;
            NN[304]=-25'd7101;
            NN[305]=-25'd2543;
            NN[306]=-25'd375;
            NN[307]=25'd136;
            NN[308]=25'd45;
            NN[309]=25'd2571;
            NN[310]=25'd9520;
            NN[311]=25'd15312;
            NN[312]=25'd20236;
            NN[313]=25'd10839;
            NN[314]=25'd2633;
            NN[315]=25'd4567;
            NN[316]=-25'd1491;
            NN[317]=25'd7322;
            NN[318]=25'd10856;
            NN[319]=25'd5887;
            NN[320]=-25'd686;
            NN[321]=25'd3960;
            NN[322]=25'd14885;
            NN[323]=25'd31993;
            NN[324]=25'd41466;
            NN[325]=25'd32967;
            NN[326]=25'd29454;
            NN[327]=25'd20317;
            NN[328]=25'd17639;
            NN[329]=25'd17484;
            NN[330]=25'd6023;
            NN[331]=-25'd7246;
            NN[332]=-25'd5595;
            NN[333]=-25'd1928;
            NN[334]=-25'd608;
            NN[335]=-25'd16;
            NN[336]=25'd97;
            NN[337]=25'd2659;
            NN[338]=25'd9794;
            NN[339]=25'd16255;
            NN[340]=25'd19715;
            NN[341]=25'd11312;
            NN[342]=25'd3626;
            NN[343]=25'd11105;
            NN[344]=25'd12158;
            NN[345]=25'd3251;
            NN[346]=-25'd5514;
            NN[347]=-25'd14955;
            NN[348]=-25'd34754;
            NN[349]=-25'd41124;
            NN[350]=-25'd17931;
            NN[351]=25'd17029;
            NN[352]=25'd35607;
            NN[353]=25'd29380;
            NN[354]=25'd23314;
            NN[355]=25'd7248;
            NN[356]=25'd7907;
            NN[357]=25'd7900;
            NN[358]=25'd390;
            NN[359]=-25'd6174;
            NN[360]=-25'd3932;
            NN[361]=25'd392;
            NN[362]=25'd379;
            NN[363]=25'd249;
            NN[364]=25'd0;
            NN[365]=25'd1369;
            NN[366]=25'd6154;
            NN[367]=25'd11858;
            NN[368]=25'd12749;
            NN[369]=25'd5951;
            NN[370]=25'd3440;
            NN[371]=25'd4048;
            NN[372]=25'd627;
            NN[373]=-25'd8836;
            NN[374]=-25'd18884;
            NN[375]=-25'd42754;
            NN[376]=-25'd64752;
            NN[377]=-25'd67022;
            NN[378]=-25'd30363;
            NN[379]=25'd4879;
            NN[380]=25'd17291;
            NN[381]=25'd14275;
            NN[382]=25'd14495;
            NN[383]=25'd7361;
            NN[384]=25'd10104;
            NN[385]=25'd5142;
            NN[386]=-25'd335;
            NN[387]=-25'd1466;
            NN[388]=25'd3;
            NN[389]=25'd709;
            NN[390]=-25'd93;
            NN[391]=-25'd107;
        end
        15:begin
            NN[0]=-25'd3;
            NN[1]=25'd639;
            NN[2]=25'd3115;
            NN[3]=25'd6102;
            NN[4]=25'd5115;
            NN[5]=25'd2601;
            NN[6]=-25'd2066;
            NN[7]=-25'd4343;
            NN[8]=-25'd11010;
            NN[9]=-25'd22533;
            NN[10]=-25'd32146;
            NN[11]=-25'd51265;
            NN[12]=-25'd65505;
            NN[13]=-25'd57504;
            NN[14]=-25'd24149;
            NN[15]=-25'd2408;
            NN[16]=25'd5394;
            NN[17]=25'd18274;
            NN[18]=25'd32837;
            NN[19]=25'd32442;
            NN[20]=25'd20354;
            NN[21]=25'd13331;
            NN[22]=25'd12893;
            NN[23]=25'd8419;
            NN[24]=25'd1733;
            NN[25]=25'd545;
            NN[26]=-25'd150;
            NN[27]=-25'd3;
            NN[28]=25'd2;
            NN[29]=-25'd18;
            NN[30]=25'd910;
            NN[31]=25'd2332;
            NN[32]=25'd621;
            NN[33]=-25'd5298;
            NN[34]=-25'd6347;
            NN[35]=-25'd10945;
            NN[36]=-25'd22099;
            NN[37]=-25'd27236;
            NN[38]=-25'd31708;
            NN[39]=-25'd43560;
            NN[40]=-25'd51703;
            NN[41]=-25'd37479;
            NN[42]=-25'd18410;
            NN[43]=25'd2184;
            NN[44]=25'd4253;
            NN[45]=25'd33898;
            NN[46]=25'd41977;
            NN[47]=25'd31832;
            NN[48]=25'd29234;
            NN[49]=25'd23195;
            NN[50]=25'd18004;
            NN[51]=25'd5841;
            NN[52]=25'd187;
            NN[53]=-25'd1385;
            NN[54]=-25'd301;
            NN[55]=-25'd19;
            NN[56]=25'd18;
            NN[57]=-25'd63;
            NN[58]=25'd33;
            NN[59]=-25'd626;
            NN[60]=-25'd274;
            NN[61]=-25'd5602;
            NN[62]=-25'd6836;
            NN[63]=-25'd7809;
            NN[64]=-25'd18318;
            NN[65]=-25'd21544;
            NN[66]=-25'd30595;
            NN[67]=-25'd35887;
            NN[68]=-25'd26021;
            NN[69]=-25'd16971;
            NN[70]=-25'd9667;
            NN[71]=25'd8518;
            NN[72]=25'd11693;
            NN[73]=25'd27643;
            NN[74]=25'd23126;
            NN[75]=25'd22434;
            NN[76]=25'd17352;
            NN[77]=25'd14002;
            NN[78]=25'd4147;
            NN[79]=-25'd2415;
            NN[80]=-25'd2556;
            NN[81]=-25'd2304;
            NN[82]=-25'd256;
            NN[83]=-25'd12;
            NN[84]=25'd0;
            NN[85]=-25'd5;
            NN[86]=-25'd121;
            NN[87]=-25'd1026;
            NN[88]=-25'd758;
            NN[89]=-25'd5654;
            NN[90]=-25'd12627;
            NN[91]=-25'd18695;
            NN[92]=-25'd21748;
            NN[93]=-25'd22563;
            NN[94]=-25'd30328;
            NN[95]=-25'd24224;
            NN[96]=-25'd12910;
            NN[97]=25'd1621;
            NN[98]=25'd6451;
            NN[99]=25'd5924;
            NN[100]=25'd1815;
            NN[101]=25'd7323;
            NN[102]=25'd7487;
            NN[103]=25'd1696;
            NN[104]=-25'd217;
            NN[105]=-25'd3598;
            NN[106]=-25'd4378;
            NN[107]=-25'd5834;
            NN[108]=-25'd2507;
            NN[109]=-25'd885;
            NN[110]=25'd204;
            NN[111]=-25'd29;
            NN[112]=25'd110;
            NN[113]=25'd0;
            NN[114]=25'd144;
            NN[115]=-25'd505;
            NN[116]=-25'd3395;
            NN[117]=-25'd10203;
            NN[118]=-25'd20250;
            NN[119]=-25'd23823;
            NN[120]=-25'd27578;
            NN[121]=-25'd29586;
            NN[122]=-25'd29434;
            NN[123]=-25'd18396;
            NN[124]=-25'd10121;
            NN[125]=25'd5109;
            NN[126]=25'd6221;
            NN[127]=-25'd2462;
            NN[128]=-25'd10130;
            NN[129]=-25'd8733;
            NN[130]=-25'd9465;
            NN[131]=-25'd10084;
            NN[132]=-25'd12466;
            NN[133]=-25'd15193;
            NN[134]=-25'd13033;
            NN[135]=-25'd11910;
            NN[136]=-25'd7041;
            NN[137]=-25'd1164;
            NN[138]=25'd325;
            NN[139]=25'd0;
            NN[140]=25'd0;
            NN[141]=25'd320;
            NN[142]=25'd140;
            NN[143]=-25'd1385;
            NN[144]=-25'd3645;
            NN[145]=-25'd12619;
            NN[146]=-25'd21000;
            NN[147]=-25'd26830;
            NN[148]=-25'd26378;
            NN[149]=-25'd25560;
            NN[150]=-25'd23606;
            NN[151]=-25'd15870;
            NN[152]=-25'd4497;
            NN[153]=25'd4324;
            NN[154]=25'd9001;
            NN[155]=-25'd6648;
            NN[156]=-25'd20426;
            NN[157]=-25'd20558;
            NN[158]=-25'd21125;
            NN[159]=-25'd17422;
            NN[160]=-25'd24925;
            NN[161]=-25'd26961;
            NN[162]=-25'd20292;
            NN[163]=-25'd12469;
            NN[164]=-25'd4103;
            NN[165]=-25'd916;
            NN[166]=-25'd135;
            NN[167]=25'd0;
            NN[168]=25'd0;
            NN[169]=-25'd4;
            NN[170]=-25'd302;
            NN[171]=-25'd2443;
            NN[172]=-25'd6557;
            NN[173]=-25'd13249;
            NN[174]=-25'd22010;
            NN[175]=-25'd26462;
            NN[176]=-25'd24637;
            NN[177]=-25'd24397;
            NN[178]=-25'd20668;
            NN[179]=-25'd15632;
            NN[180]=-25'd3012;
            NN[181]=25'd2292;
            NN[182]=25'd1876;
            NN[183]=-25'd12008;
            NN[184]=-25'd22548;
            NN[185]=-25'd27269;
            NN[186]=-25'd30518;
            NN[187]=-25'd26708;
            NN[188]=-25'd32501;
            NN[189]=-25'd28330;
            NN[190]=-25'd20123;
            NN[191]=-25'd10107;
            NN[192]=-25'd2459;
            NN[193]=-25'd621;
            NN[194]=-25'd97;
            NN[195]=25'd0;
            NN[196]=25'd0;
            NN[197]=-25'd3;
            NN[198]=-25'd828;
            NN[199]=-25'd2861;
            NN[200]=-25'd6488;
            NN[201]=-25'd10861;
            NN[202]=-25'd16450;
            NN[203]=-25'd19764;
            NN[204]=-25'd17042;
            NN[205]=-25'd20191;
            NN[206]=-25'd18021;
            NN[207]=-25'd12118;
            NN[208]=-25'd7397;
            NN[209]=-25'd8327;
            NN[210]=-25'd10175;
            NN[211]=-25'd14194;
            NN[212]=-25'd17214;
            NN[213]=-25'd23908;
            NN[214]=-25'd26020;
            NN[215]=-25'd27202;
            NN[216]=-25'd28396;
            NN[217]=-25'd24313;
            NN[218]=-25'd16315;
            NN[219]=-25'd8267;
            NN[220]=-25'd2401;
            NN[221]=-25'd656;
            NN[222]=-25'd50;
            NN[223]=25'd0;
            NN[224]=25'd0;
            NN[225]=25'd0;
            NN[226]=-25'd937;
            NN[227]=-25'd2374;
            NN[228]=-25'd3848;
            NN[229]=-25'd2374;
            NN[230]=-25'd5226;
            NN[231]=-25'd1102;
            NN[232]=-25'd4498;
            NN[233]=-25'd10566;
            NN[234]=-25'd9084;
            NN[235]=-25'd13176;
            NN[236]=-25'd12635;
            NN[237]=-25'd15056;
            NN[238]=-25'd7439;
            NN[239]=-25'd6779;
            NN[240]=-25'd11358;
            NN[241]=-25'd15267;
            NN[242]=-25'd19926;
            NN[243]=-25'd20769;
            NN[244]=-25'd24659;
            NN[245]=-25'd20438;
            NN[246]=-25'd11267;
            NN[247]=-25'd6887;
            NN[248]=-25'd1750;
            NN[249]=-25'd794;
            NN[250]=-25'd7;
            NN[251]=25'd0;
            NN[252]=25'd0;
            NN[253]=25'd0;
            NN[254]=-25'd733;
            NN[255]=-25'd1584;
            NN[256]=25'd1942;
            NN[257]=25'd5490;
            NN[258]=25'd10632;
            NN[259]=25'd15097;
            NN[260]=25'd772;
            NN[261]=-25'd282;
            NN[262]=-25'd965;
            NN[263]=-25'd8400;
            NN[264]=-25'd8338;
            NN[265]=-25'd6091;
            NN[266]=-25'd254;
            NN[267]=25'd2500;
            NN[268]=-25'd3953;
            NN[269]=-25'd5670;
            NN[270]=-25'd11779;
            NN[271]=-25'd16955;
            NN[272]=-25'd20689;
            NN[273]=-25'd16347;
            NN[274]=-25'd8950;
            NN[275]=-25'd6814;
            NN[276]=-25'd2481;
            NN[277]=-25'd893;
            NN[278]=-25'd4;
            NN[279]=25'd0;
            NN[280]=25'd0;
            NN[281]=25'd0;
            NN[282]=-25'd248;
            NN[283]=25'd475;
            NN[284]=25'd5863;
            NN[285]=25'd13440;
            NN[286]=25'd18080;
            NN[287]=25'd21000;
            NN[288]=25'd18201;
            NN[289]=25'd13302;
            NN[290]=25'd13974;
            NN[291]=25'd10511;
            NN[292]=25'd13774;
            NN[293]=25'd16318;
            NN[294]=25'd13611;
            NN[295]=25'd14317;
            NN[296]=25'd7629;
            NN[297]=25'd4317;
            NN[298]=-25'd2944;
            NN[299]=-25'd7984;
            NN[300]=-25'd11377;
            NN[301]=-25'd9999;
            NN[302]=-25'd6962;
            NN[303]=-25'd6121;
            NN[304]=-25'd2642;
            NN[305]=-25'd1089;
            NN[306]=25'd0;
            NN[307]=25'd0;
            NN[308]=25'd0;
            NN[309]=25'd0;
            NN[310]=-25'd72;
            NN[311]=25'd567;
            NN[312]=25'd4414;
            NN[313]=25'd6422;
            NN[314]=25'd8514;
            NN[315]=25'd14353;
            NN[316]=25'd22232;
            NN[317]=25'd24113;
            NN[318]=25'd20327;
            NN[319]=25'd25539;
            NN[320]=25'd27296;
            NN[321]=25'd28293;
            NN[322]=25'd24948;
            NN[323]=25'd26374;
            NN[324]=25'd20070;
            NN[325]=25'd15952;
            NN[326]=25'd11691;
            NN[327]=25'd1804;
            NN[328]=-25'd5656;
            NN[329]=-25'd4534;
            NN[330]=-25'd1943;
            NN[331]=-25'd1816;
            NN[332]=-25'd196;
            NN[333]=-25'd9;
            NN[334]=25'd0;
            NN[335]=25'd0;
            NN[336]=25'd0;
            NN[337]=25'd0;
            NN[338]=25'd0;
            NN[339]=25'd0;
            NN[340]=-25'd161;
            NN[341]=-25'd725;
            NN[342]=25'd30;
            NN[343]=25'd2873;
            NN[344]=25'd5826;
            NN[345]=25'd8268;
            NN[346]=25'd9868;
            NN[347]=25'd11307;
            NN[348]=25'd10202;
            NN[349]=25'd16039;
            NN[350]=25'd18326;
            NN[351]=25'd19866;
            NN[352]=25'd17394;
            NN[353]=25'd15280;
            NN[354]=25'd11872;
            NN[355]=25'd4329;
            NN[356]=-25'd976;
            NN[357]=-25'd833;
            NN[358]=25'd783;
            NN[359]=-25'd165;
            NN[360]=-25'd1;
            NN[361]=25'd0;
            NN[362]=25'd0;
            NN[363]=25'd0;
            NN[364]=25'd0;
            NN[365]=25'd0;
            NN[366]=25'd0;
            NN[367]=25'd0;
            NN[368]=25'd2;
            NN[369]=25'd11;
            NN[370]=25'd31;
            NN[371]=25'd274;
            NN[372]=25'd779;
            NN[373]=25'd737;
            NN[374]=25'd1284;
            NN[375]=25'd1699;
            NN[376]=25'd2105;
            NN[377]=25'd3621;
            NN[378]=25'd3931;
            NN[379]=25'd4460;
            NN[380]=25'd4537;
            NN[381]=25'd4962;
            NN[382]=25'd5004;
            NN[383]=25'd2734;
            NN[384]=25'd729;
            NN[385]=25'd13;
            NN[386]=25'd650;
            NN[387]=25'd244;
            NN[388]=25'd0;
            NN[389]=25'd0;
            NN[390]=25'd0;
            NN[391]=25'd0;
        end
        16:begin
            NN[0]=25'd0;
            NN[1]=25'd0;
            NN[2]=25'd0;
            NN[3]=25'd0;
            NN[4]=25'd0;
            NN[5]=25'd0;
            NN[6]=25'd0;
            NN[7]=25'd0;
            NN[8]=25'd0;
            NN[9]=25'd0;
            NN[10]=25'd0;
            NN[11]=25'd0;
            NN[12]=-25'd6;
            NN[13]=-25'd13;
            NN[14]=25'd0;
            NN[15]=25'd0;
            NN[16]=25'd0;
            NN[17]=25'd0;
            NN[18]=25'd0;
            NN[19]=25'd0;
            NN[20]=25'd0;
            NN[21]=25'd0;
            NN[22]=25'd0;
            NN[23]=25'd0;
            NN[24]=25'd0;
            NN[25]=25'd0;
            NN[26]=25'd0;
            NN[27]=25'd0;
            NN[28]=25'd0;
            NN[29]=25'd0;
            NN[30]=25'd0;
            NN[31]=25'd0;
            NN[32]=25'd0;
            NN[33]=25'd0;
            NN[34]=25'd0;
            NN[35]=-25'd1;
            NN[36]=-25'd23;
            NN[37]=-25'd69;
            NN[38]=-25'd169;
            NN[39]=-25'd122;
            NN[40]=-25'd95;
            NN[41]=-25'd86;
            NN[42]=-25'd93;
            NN[43]=-25'd97;
            NN[44]=-25'd188;
            NN[45]=-25'd122;
            NN[46]=-25'd67;
            NN[47]=-25'd45;
            NN[48]=-25'd35;
            NN[49]=-25'd37;
            NN[50]=-25'd4;
            NN[51]=25'd0;
            NN[52]=25'd0;
            NN[53]=25'd0;
            NN[54]=25'd0;
            NN[55]=25'd0;
            NN[56]=25'd0;
            NN[57]=25'd0;
            NN[58]=25'd0;
            NN[59]=25'd0;
            NN[60]=-25'd1;
            NN[61]=25'd0;
            NN[62]=-25'd7;
            NN[63]=-25'd43;
            NN[64]=-25'd144;
            NN[65]=-25'd561;
            NN[66]=-25'd946;
            NN[67]=-25'd1154;
            NN[68]=-25'd1588;
            NN[69]=-25'd2081;
            NN[70]=-25'd2349;
            NN[71]=-25'd2480;
            NN[72]=-25'd2503;
            NN[73]=-25'd1972;
            NN[74]=-25'd1091;
            NN[75]=-25'd1329;
            NN[76]=-25'd611;
            NN[77]=-25'd532;
            NN[78]=-25'd406;
            NN[79]=-25'd118;
            NN[80]=-25'd61;
            NN[81]=-25'd25;
            NN[82]=25'd0;
            NN[83]=25'd0;
            NN[84]=25'd0;
            NN[85]=25'd0;
            NN[86]=-25'd2;
            NN[87]=-25'd6;
            NN[88]=-25'd9;
            NN[89]=-25'd79;
            NN[90]=-25'd189;
            NN[91]=-25'd590;
            NN[92]=-25'd1099;
            NN[93]=-25'd1902;
            NN[94]=-25'd3064;
            NN[95]=-25'd4779;
            NN[96]=-25'd5830;
            NN[97]=-25'd6822;
            NN[98]=-25'd9343;
            NN[99]=-25'd9818;
            NN[100]=-25'd9889;
            NN[101]=-25'd9000;
            NN[102]=-25'd5697;
            NN[103]=-25'd6110;
            NN[104]=-25'd3202;
            NN[105]=-25'd843;
            NN[106]=25'd107;
            NN[107]=25'd810;
            NN[108]=25'd50;
            NN[109]=-25'd27;
            NN[110]=-25'd46;
            NN[111]=25'd0;
            NN[112]=25'd0;
            NN[113]=25'd0;
            NN[114]=25'd5;
            NN[115]=-25'd28;
            NN[116]=-25'd163;
            NN[117]=-25'd927;
            NN[118]=-25'd2220;
            NN[119]=-25'd3002;
            NN[120]=-25'd2510;
            NN[121]=-25'd1673;
            NN[122]=-25'd695;
            NN[123]=25'd1061;
            NN[124]=25'd9205;
            NN[125]=25'd9537;
            NN[126]=25'd15104;
            NN[127]=25'd11730;
            NN[128]=25'd3873;
            NN[129]=-25'd4012;
            NN[130]=-25'd6066;
            NN[131]=-25'd5658;
            NN[132]=-25'd1945;
            NN[133]=-25'd5795;
            NN[134]=-25'd6729;
            NN[135]=-25'd5577;
            NN[136]=-25'd714;
            NN[137]=25'd581;
            NN[138]=25'd353;
            NN[139]=25'd19;
            NN[140]=25'd0;
            NN[141]=25'd0;
            NN[142]=-25'd15;
            NN[143]=-25'd441;
            NN[144]=-25'd1159;
            NN[145]=-25'd2840;
            NN[146]=-25'd4794;
            NN[147]=-25'd4410;
            NN[148]=-25'd4339;
            NN[149]=-25'd597;
            NN[150]=-25'd2924;
            NN[151]=25'd7704;
            NN[152]=25'd17586;
            NN[153]=25'd17213;
            NN[154]=25'd18895;
            NN[155]=25'd16974;
            NN[156]=25'd16199;
            NN[157]=25'd17706;
            NN[158]=25'd4869;
            NN[159]=25'd5690;
            NN[160]=25'd3446;
            NN[161]=-25'd2343;
            NN[162]=-25'd9085;
            NN[163]=-25'd10018;
            NN[164]=-25'd2714;
            NN[165]=25'd1742;
            NN[166]=-25'd6;
            NN[167]=-25'd120;
            NN[168]=25'd0;
            NN[169]=25'd0;
            NN[170]=-25'd73;
            NN[171]=-25'd1152;
            NN[172]=-25'd2119;
            NN[173]=-25'd3803;
            NN[174]=-25'd6436;
            NN[175]=-25'd4769;
            NN[176]=25'd729;
            NN[177]=25'd2064;
            NN[178]=-25'd179;
            NN[179]=25'd6640;
            NN[180]=25'd11720;
            NN[181]=25'd5246;
            NN[182]=25'd7301;
            NN[183]=25'd18811;
            NN[184]=25'd12276;
            NN[185]=25'd8479;
            NN[186]=-25'd2390;
            NN[187]=25'd9311;
            NN[188]=25'd4077;
            NN[189]=-25'd505;
            NN[190]=-25'd2185;
            NN[191]=25'd4580;
            NN[192]=25'd3171;
            NN[193]=25'd2534;
            NN[194]=-25'd94;
            NN[195]=-25'd143;
            NN[196]=25'd0;
            NN[197]=-25'd52;
            NN[198]=-25'd231;
            NN[199]=-25'd1300;
            NN[200]=-25'd1573;
            NN[201]=-25'd2882;
            NN[202]=-25'd2149;
            NN[203]=25'd2582;
            NN[204]=25'd6907;
            NN[205]=25'd3306;
            NN[206]=25'd5928;
            NN[207]=-25'd3588;
            NN[208]=-25'd1229;
            NN[209]=-25'd429;
            NN[210]=-25'd10404;
            NN[211]=25'd4136;
            NN[212]=25'd3953;
            NN[213]=-25'd3544;
            NN[214]=25'd4653;
            NN[215]=-25'd1312;
            NN[216]=25'd2071;
            NN[217]=25'd7652;
            NN[218]=25'd7488;
            NN[219]=25'd17972;
            NN[220]=25'd14302;
            NN[221]=25'd1019;
            NN[222]=-25'd491;
            NN[223]=-25'd184;
            NN[224]=25'd0;
            NN[225]=-25'd68;
            NN[226]=-25'd487;
            NN[227]=-25'd1073;
            NN[228]=25'd913;
            NN[229]=25'd2860;
            NN[230]=25'd7889;
            NN[231]=25'd10370;
            NN[232]=25'd6818;
            NN[233]=25'd11809;
            NN[234]=25'd7606;
            NN[235]=25'd3603;
            NN[236]=25'd13728;
            NN[237]=25'd11059;
            NN[238]=-25'd12458;
            NN[239]=-25'd10007;
            NN[240]=25'd3763;
            NN[241]=-25'd2109;
            NN[242]=25'd9473;
            NN[243]=25'd9282;
            NN[244]=25'd4136;
            NN[245]=25'd10352;
            NN[246]=25'd18186;
            NN[247]=25'd20675;
            NN[248]=25'd16135;
            NN[249]=25'd2813;
            NN[250]=25'd828;
            NN[251]=25'd63;
            NN[252]=-25'd1;
            NN[253]=-25'd51;
            NN[254]=-25'd965;
            NN[255]=-25'd1423;
            NN[256]=25'd1580;
            NN[257]=25'd7299;
            NN[258]=25'd12554;
            NN[259]=25'd12516;
            NN[260]=25'd15192;
            NN[261]=25'd15321;
            NN[262]=25'd13720;
            NN[263]=25'd13439;
            NN[264]=25'd9895;
            NN[265]=-25'd149;
            NN[266]=-25'd18107;
            NN[267]=-25'd27807;
            NN[268]=-25'd18309;
            NN[269]=-25'd6167;
            NN[270]=25'd5309;
            NN[271]=25'd6948;
            NN[272]=25'd5423;
            NN[273]=25'd10529;
            NN[274]=25'd18089;
            NN[275]=25'd17630;
            NN[276]=25'd6155;
            NN[277]=25'd194;
            NN[278]=25'd2254;
            NN[279]=-25'd693;
            NN[280]=-25'd2;
            NN[281]=-25'd34;
            NN[282]=-25'd804;
            NN[283]=-25'd2636;
            NN[284]=25'd4468;
            NN[285]=25'd7573;
            NN[286]=25'd15445;
            NN[287]=25'd20022;
            NN[288]=25'd20340;
            NN[289]=25'd20343;
            NN[290]=25'd21939;
            NN[291]=25'd16155;
            NN[292]=25'd14396;
            NN[293]=25'd3607;
            NN[294]=-25'd6769;
            NN[295]=-25'd21778;
            NN[296]=-25'd27204;
            NN[297]=-25'd14575;
            NN[298]=25'd4276;
            NN[299]=25'd5425;
            NN[300]=25'd1430;
            NN[301]=25'd10526;
            NN[302]=25'd17254;
            NN[303]=25'd16318;
            NN[304]=25'd2376;
            NN[305]=-25'd3535;
            NN[306]=25'd5;
            NN[307]=25'd339;
            NN[308]=-25'd1;
            NN[309]=-25'd67;
            NN[310]=-25'd550;
            NN[311]=-25'd1807;
            NN[312]=25'd2097;
            NN[313]=25'd10494;
            NN[314]=25'd18927;
            NN[315]=25'd28026;
            NN[316]=25'd22436;
            NN[317]=25'd24840;
            NN[318]=25'd16602;
            NN[319]=25'd10674;
            NN[320]=25'd15699;
            NN[321]=25'd24850;
            NN[322]=25'd27078;
            NN[323]=-25'd2584;
            NN[324]=-25'd17878;
            NN[325]=-25'd12806;
            NN[326]=-25'd6496;
            NN[327]=-25'd499;
            NN[328]=25'd4941;
            NN[329]=25'd15695;
            NN[330]=25'd23630;
            NN[331]=25'd21760;
            NN[332]=25'd14247;
            NN[333]=25'd3014;
            NN[334]=25'd1921;
            NN[335]=25'd238;
            NN[336]=-25'd1;
            NN[337]=-25'd43;
            NN[338]=-25'd328;
            NN[339]=-25'd40;
            NN[340]=25'd311;
            NN[341]=25'd8439;
            NN[342]=25'd11622;
            NN[343]=25'd14436;
            NN[344]=25'd8242;
            NN[345]=25'd11437;
            NN[346]=-25'd2504;
            NN[347]=-25'd1337;
            NN[348]=25'd16929;
            NN[349]=25'd35538;
            NN[350]=25'd24614;
            NN[351]=25'd4016;
            NN[352]=-25'd1533;
            NN[353]=-25'd3906;
            NN[354]=-25'd5210;
            NN[355]=25'd7982;
            NN[356]=25'd15913;
            NN[357]=25'd24602;
            NN[358]=25'd20906;
            NN[359]=25'd20388;
            NN[360]=25'd13609;
            NN[361]=25'd2891;
            NN[362]=25'd248;
            NN[363]=-25'd126;
            NN[364]=25'd0;
            NN[365]=-25'd9;
            NN[366]=-25'd100;
            NN[367]=-25'd61;
            NN[368]=-25'd2795;
            NN[369]=-25'd1606;
            NN[370]=-25'd2998;
            NN[371]=-25'd4504;
            NN[372]=-25'd8651;
            NN[373]=-25'd6261;
            NN[374]=-25'd12174;
            NN[375]=25'd5771;
            NN[376]=25'd24548;
            NN[377]=25'd33198;
            NN[378]=25'd11382;
            NN[379]=25'd16852;
            NN[380]=25'd5124;
            NN[381]=-25'd7066;
            NN[382]=25'd2391;
            NN[383]=25'd6356;
            NN[384]=25'd8826;
            NN[385]=25'd1120;
            NN[386]=25'd2903;
            NN[387]=25'd5470;
            NN[388]=25'd2172;
            NN[389]=25'd291;
            NN[390]=-25'd551;
            NN[391]=-25'd135;
        end
        17:begin
            NN[0]=-25'd12;
            NN[1]=-25'd53;
            NN[2]=-25'd64;
            NN[3]=-25'd916;
            NN[4]=-25'd5078;
            NN[5]=-25'd8517;
            NN[6]=-25'd16501;
            NN[7]=-25'd24963;
            NN[8]=-25'd25437;
            NN[9]=-25'd24165;
            NN[10]=-25'd11461;
            NN[11]=25'd12388;
            NN[12]=25'd26992;
            NN[13]=25'd36377;
            NN[14]=25'd22123;
            NN[15]=25'd13722;
            NN[16]=-25'd2947;
            NN[17]=-25'd1305;
            NN[18]=-25'd4952;
            NN[19]=-25'd7491;
            NN[20]=-25'd15876;
            NN[21]=-25'd17428;
            NN[22]=-25'd15749;
            NN[23]=-25'd11240;
            NN[24]=-25'd5429;
            NN[25]=-25'd131;
            NN[26]=-25'd425;
            NN[27]=-25'd29;
            NN[28]=-25'd4;
            NN[29]=-25'd115;
            NN[30]=-25'd134;
            NN[31]=-25'd882;
            NN[32]=-25'd5105;
            NN[33]=-25'd13456;
            NN[34]=-25'd20641;
            NN[35]=-25'd23517;
            NN[36]=-25'd18516;
            NN[37]=-25'd10171;
            NN[38]=-25'd8484;
            NN[39]=25'd2668;
            NN[40]=25'd23175;
            NN[41]=25'd34074;
            NN[42]=25'd24931;
            NN[43]=25'd8459;
            NN[44]=-25'd562;
            NN[45]=-25'd11402;
            NN[46]=-25'd13922;
            NN[47]=-25'd20342;
            NN[48]=-25'd27007;
            NN[49]=-25'd25599;
            NN[50]=-25'd18429;
            NN[51]=-25'd13510;
            NN[52]=-25'd8608;
            NN[53]=-25'd1356;
            NN[54]=-25'd969;
            NN[55]=-25'd133;
            NN[56]=25'd0;
            NN[57]=-25'd58;
            NN[58]=-25'd310;
            NN[59]=-25'd834;
            NN[60]=-25'd6780;
            NN[61]=-25'd15897;
            NN[62]=-25'd17684;
            NN[63]=-25'd9585;
            NN[64]=25'd3051;
            NN[65]=25'd7686;
            NN[66]=25'd2623;
            NN[67]=25'd7220;
            NN[68]=25'd31615;
            NN[69]=25'd19242;
            NN[70]=25'd4521;
            NN[71]=25'd4254;
            NN[72]=25'd1779;
            NN[73]=-25'd9566;
            NN[74]=-25'd22263;
            NN[75]=-25'd26242;
            NN[76]=-25'd25641;
            NN[77]=-25'd27322;
            NN[78]=-25'd20630;
            NN[79]=-25'd9653;
            NN[80]=-25'd8175;
            NN[81]=-25'd4317;
            NN[82]=-25'd1669;
            NN[83]=-25'd106;
            NN[84]=25'd0;
            NN[85]=-25'd39;
            NN[86]=-25'd381;
            NN[87]=-25'd2043;
            NN[88]=-25'd8501;
            NN[89]=-25'd15878;
            NN[90]=-25'd13767;
            NN[91]=25'd396;
            NN[92]=25'd15417;
            NN[93]=25'd22236;
            NN[94]=25'd7755;
            NN[95]=25'd21718;
            NN[96]=25'd34147;
            NN[97]=25'd15186;
            NN[98]=-25'd1994;
            NN[99]=-25'd6529;
            NN[100]=25'd1197;
            NN[101]=-25'd12881;
            NN[102]=-25'd19458;
            NN[103]=-25'd10488;
            NN[104]=-25'd10280;
            NN[105]=-25'd14407;
            NN[106]=-25'd14297;
            NN[107]=-25'd4769;
            NN[108]=-25'd4434;
            NN[109]=-25'd6176;
            NN[110]=-25'd1426;
            NN[111]=-25'd27;
            NN[112]=-25'd9;
            NN[113]=-25'd4;
            NN[114]=-25'd288;
            NN[115]=-25'd3990;
            NN[116]=-25'd11826;
            NN[117]=-25'd11495;
            NN[118]=-25'd4653;
            NN[119]=25'd5353;
            NN[120]=25'd14335;
            NN[121]=25'd21653;
            NN[122]=25'd21707;
            NN[123]=25'd24168;
            NN[124]=25'd19275;
            NN[125]=25'd1731;
            NN[126]=-25'd12179;
            NN[127]=-25'd6054;
            NN[128]=-25'd11046;
            NN[129]=-25'd10852;
            NN[130]=-25'd3427;
            NN[131]=25'd107;
            NN[132]=-25'd590;
            NN[133]=-25'd8836;
            NN[134]=-25'd4570;
            NN[135]=-25'd1551;
            NN[136]=-25'd4261;
            NN[137]=-25'd4708;
            NN[138]=-25'd598;
            NN[139]=-25'd14;
            NN[140]=25'd0;
            NN[141]=-25'd27;
            NN[142]=-25'd371;
            NN[143]=-25'd5747;
            NN[144]=-25'd11996;
            NN[145]=-25'd4883;
            NN[146]=25'd3800;
            NN[147]=25'd9000;
            NN[148]=25'd9809;
            NN[149]=25'd15166;
            NN[150]=25'd12463;
            NN[151]=-25'd2240;
            NN[152]=-25'd260;
            NN[153]=-25'd12621;
            NN[154]=-25'd15084;
            NN[155]=-25'd5443;
            NN[156]=-25'd7396;
            NN[157]=-25'd4058;
            NN[158]=25'd3835;
            NN[159]=25'd4391;
            NN[160]=25'd3919;
            NN[161]=-25'd88;
            NN[162]=25'd5232;
            NN[163]=25'd3104;
            NN[164]=-25'd3900;
            NN[165]=-25'd3479;
            NN[166]=-25'd655;
            NN[167]=-25'd7;
            NN[168]=25'd0;
            NN[169]=-25'd46;
            NN[170]=-25'd515;
            NN[171]=-25'd5918;
            NN[172]=-25'd10144;
            NN[173]=-25'd6289;
            NN[174]=25'd7679;
            NN[175]=25'd18747;
            NN[176]=25'd7168;
            NN[177]=-25'd621;
            NN[178]=25'd3194;
            NN[179]=-25'd11206;
            NN[180]=-25'd1626;
            NN[181]=-25'd4329;
            NN[182]=-25'd12383;
            NN[183]=-25'd1983;
            NN[184]=-25'd11074;
            NN[185]=-25'd4362;
            NN[186]=-25'd1227;
            NN[187]=25'd1834;
            NN[188]=25'd6933;
            NN[189]=25'd9070;
            NN[190]=25'd8761;
            NN[191]=25'd1753;
            NN[192]=-25'd4563;
            NN[193]=-25'd2307;
            NN[194]=-25'd548;
            NN[195]=-25'd5;
            NN[196]=25'd0;
            NN[197]=-25'd2;
            NN[198]=-25'd565;
            NN[199]=-25'd4229;
            NN[200]=-25'd7500;
            NN[201]=-25'd6333;
            NN[202]=25'd9060;
            NN[203]=25'd17882;
            NN[204]=25'd5870;
            NN[205]=25'd4834;
            NN[206]=-25'd1143;
            NN[207]=-25'd1771;
            NN[208]=25'd110;
            NN[209]=25'd4208;
            NN[210]=-25'd556;
            NN[211]=-25'd2496;
            NN[212]=-25'd10412;
            NN[213]=-25'd6590;
            NN[214]=-25'd1767;
            NN[215]=25'd92;
            NN[216]=25'd6712;
            NN[217]=25'd6666;
            NN[218]=25'd5096;
            NN[219]=-25'd3328;
            NN[220]=-25'd5178;
            NN[221]=-25'd1589;
            NN[222]=-25'd227;
            NN[223]=25'd0;
            NN[224]=25'd0;
            NN[225]=25'd0;
            NN[226]=-25'd472;
            NN[227]=-25'd2375;
            NN[228]=-25'd7225;
            NN[229]=-25'd12222;
            NN[230]=-25'd1667;
            NN[231]=25'd8236;
            NN[232]=25'd4271;
            NN[233]=25'd459;
            NN[234]=25'd1675;
            NN[235]=25'd13026;
            NN[236]=25'd18600;
            NN[237]=25'd20784;
            NN[238]=25'd18838;
            NN[239]=25'd9431;
            NN[240]=25'd538;
            NN[241]=25'd4703;
            NN[242]=25'd5643;
            NN[243]=-25'd564;
            NN[244]=25'd1763;
            NN[245]=25'd4151;
            NN[246]=-25'd2504;
            NN[247]=-25'd3062;
            NN[248]=-25'd2588;
            NN[249]=-25'd517;
            NN[250]=-25'd117;
            NN[251]=25'd0;
            NN[252]=25'd0;
            NN[253]=25'd0;
            NN[254]=-25'd114;
            NN[255]=-25'd1297;
            NN[256]=-25'd7327;
            NN[257]=-25'd20283;
            NN[258]=-25'd22358;
            NN[259]=-25'd11546;
            NN[260]=25'd4919;
            NN[261]=25'd2593;
            NN[262]=25'd1446;
            NN[263]=25'd10053;
            NN[264]=25'd21594;
            NN[265]=25'd34691;
            NN[266]=25'd28257;
            NN[267]=25'd23579;
            NN[268]=25'd22163;
            NN[269]=25'd12054;
            NN[270]=25'd11984;
            NN[271]=25'd8766;
            NN[272]=25'd9324;
            NN[273]=25'd2010;
            NN[274]=-25'd1525;
            NN[275]=-25'd401;
            NN[276]=-25'd1364;
            NN[277]=-25'd395;
            NN[278]=-25'd266;
            NN[279]=25'd0;
            NN[280]=25'd0;
            NN[281]=25'd0;
            NN[282]=-25'd5;
            NN[283]=-25'd818;
            NN[284]=-25'd5784;
            NN[285]=-25'd15750;
            NN[286]=-25'd21707;
            NN[287]=-25'd17960;
            NN[288]=-25'd6229;
            NN[289]=-25'd3169;
            NN[290]=25'd3352;
            NN[291]=25'd10924;
            NN[292]=25'd11772;
            NN[293]=25'd9947;
            NN[294]=25'd12998;
            NN[295]=25'd19872;
            NN[296]=25'd22026;
            NN[297]=25'd9555;
            NN[298]=25'd13931;
            NN[299]=25'd14614;
            NN[300]=25'd5176;
            NN[301]=-25'd1522;
            NN[302]=-25'd2924;
            NN[303]=-25'd1638;
            NN[304]=-25'd1005;
            NN[305]=-25'd477;
            NN[306]=-25'd87;
            NN[307]=25'd0;
            NN[308]=25'd0;
            NN[309]=25'd0;
            NN[310]=-25'd3;
            NN[311]=-25'd232;
            NN[312]=-25'd3202;
            NN[313]=-25'd6415;
            NN[314]=-25'd7649;
            NN[315]=-25'd9798;
            NN[316]=-25'd13367;
            NN[317]=-25'd15087;
            NN[318]=-25'd10205;
            NN[319]=-25'd10399;
            NN[320]=-25'd11794;
            NN[321]=-25'd8069;
            NN[322]=-25'd629;
            NN[323]=25'd6112;
            NN[324]=25'd5936;
            NN[325]=25'd5488;
            NN[326]=25'd2897;
            NN[327]=25'd1474;
            NN[328]=25'd152;
            NN[329]=-25'd1212;
            NN[330]=-25'd1149;
            NN[331]=-25'd298;
            NN[332]=-25'd75;
            NN[333]=-25'd57;
            NN[334]=-25'd61;
            NN[335]=25'd0;
            NN[336]=25'd0;
            NN[337]=25'd0;
            NN[338]=25'd0;
            NN[339]=25'd0;
            NN[340]=-25'd468;
            NN[341]=-25'd1088;
            NN[342]=-25'd1555;
            NN[343]=-25'd1255;
            NN[344]=-25'd1718;
            NN[345]=-25'd3121;
            NN[346]=-25'd4693;
            NN[347]=-25'd4334;
            NN[348]=-25'd4965;
            NN[349]=-25'd5721;
            NN[350]=-25'd5550;
            NN[351]=-25'd5495;
            NN[352]=-25'd4380;
            NN[353]=-25'd2828;
            NN[354]=-25'd1997;
            NN[355]=-25'd1647;
            NN[356]=-25'd1029;
            NN[357]=-25'd538;
            NN[358]=-25'd110;
            NN[359]=-25'd13;
            NN[360]=25'd0;
            NN[361]=25'd0;
            NN[362]=25'd0;
            NN[363]=25'd0;
            NN[364]=25'd0;
            NN[365]=25'd0;
            NN[366]=25'd0;
            NN[367]=25'd0;
            NN[368]=25'd0;
            NN[369]=-25'd2;
            NN[370]=-25'd4;
            NN[371]=-25'd23;
            NN[372]=-25'd42;
            NN[373]=-25'd61;
            NN[374]=-25'd256;
            NN[375]=-25'd191;
            NN[376]=-25'd238;
            NN[377]=-25'd274;
            NN[378]=-25'd393;
            NN[379]=-25'd373;
            NN[380]=-25'd335;
            NN[381]=-25'd298;
            NN[382]=-25'd191;
            NN[383]=-25'd98;
            NN[384]=-25'd95;
            NN[385]=-25'd46;
            NN[386]=-25'd47;
            NN[387]=-25'd8;
            NN[388]=25'd0;
            NN[389]=25'd0;
            NN[390]=25'd0;
            NN[391]=25'd0;
        end
        18:begin
            NN[0]=25'd0;
            NN[1]=25'd0;
            NN[2]=25'd0;
            NN[3]=25'd0;
            NN[4]=25'd0;
            NN[5]=25'd0;
            NN[6]=25'd0;
            NN[7]=25'd0;
            NN[8]=25'd0;
            NN[9]=25'd0;
            NN[10]=25'd0;
            NN[11]=25'd0;
            NN[12]=-25'd32;
            NN[13]=-25'd71;
            NN[14]=25'd0;
            NN[15]=25'd0;
            NN[16]=25'd0;
            NN[17]=25'd0;
            NN[18]=25'd0;
            NN[19]=25'd0;
            NN[20]=25'd0;
            NN[21]=25'd0;
            NN[22]=25'd0;
            NN[23]=25'd0;
            NN[24]=25'd0;
            NN[25]=25'd0;
            NN[26]=25'd0;
            NN[27]=25'd0;
            NN[28]=25'd0;
            NN[29]=25'd0;
            NN[30]=25'd0;
            NN[31]=25'd0;
            NN[32]=25'd0;
            NN[33]=25'd0;
            NN[34]=-25'd2;
            NN[35]=-25'd7;
            NN[36]=-25'd30;
            NN[37]=-25'd97;
            NN[38]=-25'd235;
            NN[39]=-25'd266;
            NN[40]=-25'd378;
            NN[41]=-25'd215;
            NN[42]=-25'd92;
            NN[43]=-25'd305;
            NN[44]=-25'd757;
            NN[45]=-25'd409;
            NN[46]=-25'd77;
            NN[47]=-25'd69;
            NN[48]=-25'd55;
            NN[49]=-25'd18;
            NN[50]=-25'd8;
            NN[51]=-25'd3;
            NN[52]=25'd0;
            NN[53]=25'd0;
            NN[54]=25'd0;
            NN[55]=25'd0;
            NN[56]=25'd0;
            NN[57]=25'd0;
            NN[58]=25'd0;
            NN[59]=-25'd2;
            NN[60]=-25'd2;
            NN[61]=25'd0;
            NN[62]=-25'd4;
            NN[63]=-25'd53;
            NN[64]=-25'd145;
            NN[65]=-25'd412;
            NN[66]=-25'd776;
            NN[67]=-25'd952;
            NN[68]=-25'd1315;
            NN[69]=-25'd1387;
            NN[70]=-25'd1532;
            NN[71]=-25'd1703;
            NN[72]=-25'd1894;
            NN[73]=-25'd1433;
            NN[74]=-25'd974;
            NN[75]=-25'd689;
            NN[76]=-25'd373;
            NN[77]=-25'd366;
            NN[78]=-25'd246;
            NN[79]=-25'd37;
            NN[80]=-25'd2;
            NN[81]=25'd0;
            NN[82]=25'd0;
            NN[83]=25'd0;
            NN[84]=25'd0;
            NN[85]=25'd0;
            NN[86]=25'd0;
            NN[87]=-25'd9;
            NN[88]=-25'd8;
            NN[89]=-25'd22;
            NN[90]=-25'd72;
            NN[91]=-25'd196;
            NN[92]=-25'd611;
            NN[93]=-25'd1198;
            NN[94]=-25'd2128;
            NN[95]=-25'd2851;
            NN[96]=-25'd3584;
            NN[97]=-25'd4658;
            NN[98]=-25'd6140;
            NN[99]=-25'd7371;
            NN[100]=-25'd6812;
            NN[101]=-25'd4858;
            NN[102]=-25'd2905;
            NN[103]=-25'd2474;
            NN[104]=-25'd1956;
            NN[105]=-25'd1267;
            NN[106]=-25'd507;
            NN[107]=-25'd177;
            NN[108]=-25'd56;
            NN[109]=-25'd8;
            NN[110]=25'd0;
            NN[111]=25'd0;
            NN[112]=25'd0;
            NN[113]=25'd0;
            NN[114]=25'd0;
            NN[115]=-25'd8;
            NN[116]=-25'd52;
            NN[117]=-25'd284;
            NN[118]=-25'd651;
            NN[119]=-25'd1190;
            NN[120]=-25'd2274;
            NN[121]=-25'd4591;
            NN[122]=-25'd6706;
            NN[123]=-25'd9152;
            NN[124]=-25'd12397;
            NN[125]=-25'd15363;
            NN[126]=-25'd19997;
            NN[127]=-25'd23021;
            NN[128]=-25'd23152;
            NN[129]=-25'd17553;
            NN[130]=-25'd13011;
            NN[131]=-25'd10766;
            NN[132]=-25'd7668;
            NN[133]=-25'd5740;
            NN[134]=-25'd3343;
            NN[135]=-25'd1632;
            NN[136]=-25'd687;
            NN[137]=-25'd264;
            NN[138]=-25'd70;
            NN[139]=-25'd3;
            NN[140]=25'd0;
            NN[141]=25'd0;
            NN[142]=25'd0;
            NN[143]=-25'd129;
            NN[144]=-25'd379;
            NN[145]=-25'd1650;
            NN[146]=-25'd4219;
            NN[147]=-25'd6355;
            NN[148]=-25'd8857;
            NN[149]=-25'd12699;
            NN[150]=-25'd9461;
            NN[151]=-25'd3080;
            NN[152]=-25'd2581;
            NN[153]=-25'd1671;
            NN[154]=-25'd10028;
            NN[155]=-25'd16564;
            NN[156]=-25'd30356;
            NN[157]=-25'd29798;
            NN[158]=-25'd27567;
            NN[159]=-25'd23953;
            NN[160]=-25'd19940;
            NN[161]=-25'd16386;
            NN[162]=-25'd14186;
            NN[163]=-25'd9350;
            NN[164]=-25'd4637;
            NN[165]=-25'd1706;
            NN[166]=-25'd159;
            NN[167]=-25'd2;
            NN[168]=25'd0;
            NN[169]=-25'd5;
            NN[170]=-25'd104;
            NN[171]=-25'd564;
            NN[172]=-25'd2159;
            NN[173]=-25'd6704;
            NN[174]=-25'd11797;
            NN[175]=-25'd17483;
            NN[176]=-25'd19634;
            NN[177]=-25'd14958;
            NN[178]=-25'd8733;
            NN[179]=25'd2560;
            NN[180]=25'd7022;
            NN[181]=25'd20007;
            NN[182]=25'd24135;
            NN[183]=25'd16715;
            NN[184]=25'd14913;
            NN[185]=25'd11311;
            NN[186]=25'd9315;
            NN[187]=-25'd3380;
            NN[188]=-25'd9552;
            NN[189]=-25'd15403;
            NN[190]=-25'd20453;
            NN[191]=-25'd18680;
            NN[192]=-25'd11416;
            NN[193]=-25'd4384;
            NN[194]=-25'd1219;
            NN[195]=-25'd92;
            NN[196]=25'd0;
            NN[197]=-25'd187;
            NN[198]=-25'd544;
            NN[199]=-25'd2275;
            NN[200]=-25'd6961;
            NN[201]=-25'd14267;
            NN[202]=-25'd19092;
            NN[203]=-25'd23449;
            NN[204]=-25'd15881;
            NN[205]=-25'd3521;
            NN[206]=25'd1246;
            NN[207]=25'd7106;
            NN[208]=25'd18257;
            NN[209]=25'd29620;
            NN[210]=25'd43198;
            NN[211]=25'd50780;
            NN[212]=25'd47245;
            NN[213]=25'd30969;
            NN[214]=25'd17858;
            NN[215]=25'd8043;
            NN[216]=25'd2794;
            NN[217]=-25'd7573;
            NN[218]=-25'd21756;
            NN[219]=-25'd22497;
            NN[220]=-25'd15773;
            NN[221]=-25'd6114;
            NN[222]=-25'd1558;
            NN[223]=-25'd74;
            NN[224]=-25'd30;
            NN[225]=-25'd699;
            NN[226]=-25'd1819;
            NN[227]=-25'd5580;
            NN[228]=-25'd11042;
            NN[229]=-25'd15880;
            NN[230]=-25'd13460;
            NN[231]=-25'd17506;
            NN[232]=-25'd1257;
            NN[233]=-25'd2877;
            NN[234]=-25'd2088;
            NN[235]=-25'd5329;
            NN[236]=-25'd3909;
            NN[237]=25'd14421;
            NN[238]=25'd31243;
            NN[239]=25'd27716;
            NN[240]=25'd18010;
            NN[241]=25'd7681;
            NN[242]=25'd8044;
            NN[243]=-25'd113;
            NN[244]=-25'd2019;
            NN[245]=-25'd67;
            NN[246]=-25'd16537;
            NN[247]=-25'd20772;
            NN[248]=-25'd14392;
            NN[249]=-25'd6126;
            NN[250]=-25'd1395;
            NN[251]=-25'd91;
            NN[252]=-25'd41;
            NN[253]=-25'd980;
            NN[254]=-25'd2498;
            NN[255]=-25'd6266;
            NN[256]=-25'd14031;
            NN[257]=-25'd9208;
            NN[258]=25'd1522;
            NN[259]=-25'd851;
            NN[260]=25'd4159;
            NN[261]=25'd980;
            NN[262]=25'd5089;
            NN[263]=25'd4789;
            NN[264]=25'd8099;
            NN[265]=25'd6481;
            NN[266]=25'd16877;
            NN[267]=25'd15082;
            NN[268]=-25'd1001;
            NN[269]=-25'd2312;
            NN[270]=25'd2763;
            NN[271]=-25'd80;
            NN[272]=25'd160;
            NN[273]=-25'd6955;
            NN[274]=-25'd13504;
            NN[275]=-25'd18082;
            NN[276]=-25'd12874;
            NN[277]=-25'd5996;
            NN[278]=-25'd1899;
            NN[279]=-25'd111;
            NN[280]=-25'd55;
            NN[281]=-25'd1026;
            NN[282]=-25'd3083;
            NN[283]=-25'd5567;
            NN[284]=-25'd9410;
            NN[285]=25'd613;
            NN[286]=25'd12636;
            NN[287]=25'd10162;
            NN[288]=25'd15793;
            NN[289]=25'd9627;
            NN[290]=25'd14122;
            NN[291]=25'd20805;
            NN[292]=25'd12632;
            NN[293]=-25'd7022;
            NN[294]=-25'd3600;
            NN[295]=-25'd6329;
            NN[296]=-25'd5188;
            NN[297]=25'd1909;
            NN[298]=25'd5066;
            NN[299]=25'd5136;
            NN[300]=25'd8489;
            NN[301]=25'd2660;
            NN[302]=-25'd2034;
            NN[303]=-25'd8393;
            NN[304]=-25'd12184;
            NN[305]=-25'd5567;
            NN[306]=-25'd1596;
            NN[307]=-25'd240;
            NN[308]=-25'd27;
            NN[309]=-25'd1527;
            NN[310]=-25'd4539;
            NN[311]=-25'd5459;
            NN[312]=-25'd48;
            NN[313]=25'd13667;
            NN[314]=25'd21356;
            NN[315]=25'd18075;
            NN[316]=25'd29981;
            NN[317]=25'd15973;
            NN[318]=25'd18364;
            NN[319]=25'd22144;
            NN[320]=-25'd4598;
            NN[321]=-25'd11834;
            NN[322]=-25'd1593;
            NN[323]=25'd8152;
            NN[324]=25'd13409;
            NN[325]=25'd26534;
            NN[326]=25'd21950;
            NN[327]=25'd21968;
            NN[328]=25'd34141;
            NN[329]=25'd22000;
            NN[330]=25'd12998;
            NN[331]=-25'd1891;
            NN[332]=-25'd8241;
            NN[333]=-25'd3929;
            NN[334]=-25'd1068;
            NN[335]=-25'd96;
            NN[336]=-25'd86;
            NN[337]=-25'd1145;
            NN[338]=-25'd4268;
            NN[339]=-25'd3256;
            NN[340]=25'd10476;
            NN[341]=25'd22911;
            NN[342]=25'd24177;
            NN[343]=25'd18115;
            NN[344]=25'd19471;
            NN[345]=25'd20521;
            NN[346]=25'd17507;
            NN[347]=25'd7176;
            NN[348]=-25'd16599;
            NN[349]=-25'd820;
            NN[350]=25'd20236;
            NN[351]=25'd23131;
            NN[352]=25'd24773;
            NN[353]=25'd29549;
            NN[354]=25'd27501;
            NN[355]=25'd34876;
            NN[356]=25'd38607;
            NN[357]=25'd30156;
            NN[358]=25'd18403;
            NN[359]=25'd4819;
            NN[360]=-25'd6573;
            NN[361]=-25'd2997;
            NN[362]=-25'd927;
            NN[363]=-25'd33;
            NN[364]=25'd0;
            NN[365]=-25'd458;
            NN[366]=-25'd3077;
            NN[367]=-25'd1495;
            NN[368]=25'd18366;
            NN[369]=25'd25004;
            NN[370]=25'd19068;
            NN[371]=25'd17651;
            NN[372]=25'd14493;
            NN[373]=25'd7570;
            NN[374]=25'd6850;
            NN[375]=-25'd3934;
            NN[376]=-25'd12338;
            NN[377]=25'd7473;
            NN[378]=25'd22234;
            NN[379]=25'd22093;
            NN[380]=25'd34885;
            NN[381]=25'd30022;
            NN[382]=25'd24874;
            NN[383]=25'd31378;
            NN[384]=25'd30129;
            NN[385]=25'd21736;
            NN[386]=25'd6158;
            NN[387]=-25'd7422;
            NN[388]=-25'd9814;
            NN[389]=-25'd4280;
            NN[390]=-25'd1109;
            NN[391]=-25'd54;
        end
        19:begin
            NN[0]=-25'd69;
            NN[1]=-25'd191;
            NN[2]=-25'd1836;
            NN[3]=25'd391;
            NN[4]=25'd12605;
            NN[5]=25'd13791;
            NN[6]=25'd16394;
            NN[7]=25'd12856;
            NN[8]=25'd8087;
            NN[9]=25'd3292;
            NN[10]=-25'd1356;
            NN[11]=-25'd3957;
            NN[12]=-25'd7228;
            NN[13]=25'd548;
            NN[14]=25'd860;
            NN[15]=25'd16226;
            NN[16]=25'd34750;
            NN[17]=25'd29650;
            NN[18]=25'd13446;
            NN[19]=25'd9692;
            NN[20]=25'd14052;
            NN[21]=25'd2284;
            NN[22]=-25'd8931;
            NN[23]=-25'd16559;
            NN[24]=-25'd11828;
            NN[25]=-25'd3625;
            NN[26]=-25'd471;
            NN[27]=-25'd10;
            NN[28]=-25'd23;
            NN[29]=-25'd10;
            NN[30]=-25'd1286;
            NN[31]=-25'd326;
            NN[32]=25'd5883;
            NN[33]=25'd6040;
            NN[34]=25'd4524;
            NN[35]=25'd7031;
            NN[36]=25'd6464;
            NN[37]=-25'd1010;
            NN[38]=25'd626;
            NN[39]=-25'd736;
            NN[40]=-25'd4319;
            NN[41]=-25'd13115;
            NN[42]=-25'd15165;
            NN[43]=25'd11968;
            NN[44]=25'd29171;
            NN[45]=25'd28851;
            NN[46]=25'd8770;
            NN[47]=25'd2088;
            NN[48]=25'd470;
            NN[49]=-25'd12565;
            NN[50]=-25'd17649;
            NN[51]=-25'd17959;
            NN[52]=-25'd11664;
            NN[53]=-25'd3918;
            NN[54]=-25'd1265;
            NN[55]=-25'd117;
            NN[56]=-25'd2;
            NN[57]=-25'd57;
            NN[58]=-25'd879;
            NN[59]=-25'd1013;
            NN[60]=25'd2327;
            NN[61]=-25'd1210;
            NN[62]=-25'd7237;
            NN[63]=-25'd97;
            NN[64]=25'd8332;
            NN[65]=-25'd1766;
            NN[66]=25'd6281;
            NN[67]=25'd7440;
            NN[68]=-25'd5498;
            NN[69]=-25'd19511;
            NN[70]=-25'd11005;
            NN[71]=25'd6146;
            NN[72]=25'd21423;
            NN[73]=25'd16320;
            NN[74]=25'd1575;
            NN[75]=-25'd9453;
            NN[76]=-25'd14196;
            NN[77]=-25'd23318;
            NN[78]=-25'd18701;
            NN[79]=-25'd19501;
            NN[80]=-25'd12282;
            NN[81]=-25'd3887;
            NN[82]=-25'd1089;
            NN[83]=-25'd20;
            NN[84]=25'd0;
            NN[85]=-25'd8;
            NN[86]=-25'd1123;
            NN[87]=-25'd3300;
            NN[88]=-25'd6327;
            NN[89]=-25'd8798;
            NN[90]=-25'd10681;
            NN[91]=25'd177;
            NN[92]=25'd3234;
            NN[93]=25'd3430;
            NN[94]=25'd7162;
            NN[95]=25'd7114;
            NN[96]=-25'd1555;
            NN[97]=-25'd8977;
            NN[98]=-25'd4257;
            NN[99]=25'd13197;
            NN[100]=25'd7903;
            NN[101]=25'd1088;
            NN[102]=-25'd9511;
            NN[103]=-25'd12940;
            NN[104]=-25'd15298;
            NN[105]=-25'd19617;
            NN[106]=-25'd21311;
            NN[107]=-25'd20214;
            NN[108]=-25'd12356;
            NN[109]=-25'd3200;
            NN[110]=-25'd586;
            NN[111]=-25'd40;
            NN[112]=25'd15;
            NN[113]=-25'd1;
            NN[114]=-25'd735;
            NN[115]=-25'd5170;
            NN[116]=-25'd9142;
            NN[117]=-25'd13640;
            NN[118]=-25'd11302;
            NN[119]=-25'd11375;
            NN[120]=-25'd7155;
            NN[121]=-25'd2043;
            NN[122]=25'd6696;
            NN[123]=25'd3013;
            NN[124]=-25'd12015;
            NN[125]=-25'd10813;
            NN[126]=25'd4268;
            NN[127]=25'd4846;
            NN[128]=-25'd8075;
            NN[129]=-25'd9071;
            NN[130]=-25'd12198;
            NN[131]=-25'd7765;
            NN[132]=-25'd8270;
            NN[133]=-25'd16125;
            NN[134]=-25'd19360;
            NN[135]=-25'd17565;
            NN[136]=-25'd10463;
            NN[137]=-25'd2788;
            NN[138]=-25'd98;
            NN[139]=-25'd10;
            NN[140]=25'd0;
            NN[141]=-25'd260;
            NN[142]=-25'd768;
            NN[143]=-25'd4381;
            NN[144]=-25'd8258;
            NN[145]=-25'd11867;
            NN[146]=-25'd14658;
            NN[147]=-25'd16484;
            NN[148]=-25'd19463;
            NN[149]=-25'd21672;
            NN[150]=-25'd19095;
            NN[151]=-25'd23829;
            NN[152]=-25'd21351;
            NN[153]=-25'd16468;
            NN[154]=-25'd12556;
            NN[155]=-25'd14296;
            NN[156]=-25'd9734;
            NN[157]=-25'd12639;
            NN[158]=-25'd11580;
            NN[159]=-25'd3603;
            NN[160]=-25'd5557;
            NN[161]=-25'd15575;
            NN[162]=-25'd14811;
            NN[163]=-25'd10964;
            NN[164]=-25'd5196;
            NN[165]=-25'd1343;
            NN[166]=-25'd197;
            NN[167]=25'd0;
            NN[168]=25'd0;
            NN[169]=-25'd93;
            NN[170]=-25'd633;
            NN[171]=-25'd3473;
            NN[172]=-25'd5611;
            NN[173]=-25'd7173;
            NN[174]=-25'd15171;
            NN[175]=-25'd23968;
            NN[176]=-25'd23506;
            NN[177]=-25'd30583;
            NN[178]=-25'd35698;
            NN[179]=-25'd38511;
            NN[180]=-25'd34908;
            NN[181]=-25'd17990;
            NN[182]=-25'd19323;
            NN[183]=-25'd15788;
            NN[184]=-25'd9267;
            NN[185]=-25'd12378;
            NN[186]=-25'd15346;
            NN[187]=-25'd6778;
            NN[188]=-25'd9335;
            NN[189]=-25'd13560;
            NN[190]=-25'd9779;
            NN[191]=-25'd5010;
            NN[192]=-25'd710;
            NN[193]=25'd495;
            NN[194]=-25'd170;
            NN[195]=25'd0;
            NN[196]=25'd0;
            NN[197]=-25'd6;
            NN[198]=-25'd507;
            NN[199]=-25'd2633;
            NN[200]=-25'd4475;
            NN[201]=-25'd6220;
            NN[202]=-25'd12555;
            NN[203]=-25'd19238;
            NN[204]=-25'd20109;
            NN[205]=-25'd20097;
            NN[206]=-25'd23430;
            NN[207]=-25'd30112;
            NN[208]=-25'd26693;
            NN[209]=-25'd19580;
            NN[210]=-25'd20387;
            NN[211]=-25'd17399;
            NN[212]=-25'd11203;
            NN[213]=-25'd18358;
            NN[214]=-25'd18599;
            NN[215]=-25'd15287;
            NN[216]=-25'd9823;
            NN[217]=-25'd6715;
            NN[218]=-25'd4487;
            NN[219]=-25'd324;
            NN[220]=25'd2540;
            NN[221]=25'd446;
            NN[222]=-25'd146;
            NN[223]=25'd0;
            NN[224]=25'd0;
            NN[225]=25'd0;
            NN[226]=-25'd705;
            NN[227]=-25'd1643;
            NN[228]=-25'd3636;
            NN[229]=-25'd8918;
            NN[230]=-25'd11817;
            NN[231]=-25'd16617;
            NN[232]=-25'd10277;
            NN[233]=-25'd8218;
            NN[234]=-25'd6714;
            NN[235]=-25'd10110;
            NN[236]=-25'd7738;
            NN[237]=-25'd13578;
            NN[238]=-25'd10734;
            NN[239]=-25'd15806;
            NN[240]=-25'd14507;
            NN[241]=-25'd19771;
            NN[242]=-25'd19063;
            NN[243]=-25'd20394;
            NN[244]=-25'd5552;
            NN[245]=-25'd588;
            NN[246]=25'd3708;
            NN[247]=25'd6141;
            NN[248]=25'd2771;
            NN[249]=25'd681;
            NN[250]=-25'd43;
            NN[251]=25'd0;
            NN[252]=25'd0;
            NN[253]=25'd0;
            NN[254]=-25'd350;
            NN[255]=-25'd613;
            NN[256]=-25'd3552;
            NN[257]=-25'd5819;
            NN[258]=-25'd8606;
            NN[259]=-25'd8722;
            NN[260]=-25'd480;
            NN[261]=-25'd3178;
            NN[262]=-25'd47;
            NN[263]=-25'd6680;
            NN[264]=-25'd6487;
            NN[265]=-25'd12098;
            NN[266]=-25'd10547;
            NN[267]=-25'd16610;
            NN[268]=-25'd13156;
            NN[269]=-25'd13157;
            NN[270]=-25'd12018;
            NN[271]=-25'd4904;
            NN[272]=25'd4739;
            NN[273]=25'd10535;
            NN[274]=25'd12201;
            NN[275]=25'd8888;
            NN[276]=25'd2736;
            NN[277]=25'd98;
            NN[278]=-25'd71;
            NN[279]=25'd0;
            NN[280]=25'd0;
            NN[281]=25'd0;
            NN[282]=-25'd39;
            NN[283]=-25'd299;
            NN[284]=-25'd52;
            NN[285]=25'd518;
            NN[286]=25'd799;
            NN[287]=25'd4430;
            NN[288]=25'd8370;
            NN[289]=25'd5328;
            NN[290]=25'd1950;
            NN[291]=-25'd4041;
            NN[292]=-25'd7949;
            NN[293]=-25'd11976;
            NN[294]=-25'd12208;
            NN[295]=-25'd4878;
            NN[296]=-25'd839;
            NN[297]=25'd5438;
            NN[298]=25'd8397;
            NN[299]=25'd14656;
            NN[300]=25'd22769;
            NN[301]=25'd19975;
            NN[302]=25'd13955;
            NN[303]=25'd8538;
            NN[304]=25'd241;
            NN[305]=-25'd531;
            NN[306]=-25'd260;
            NN[307]=25'd0;
            NN[308]=25'd0;
            NN[309]=25'd0;
            NN[310]=25'd27;
            NN[311]=-25'd201;
            NN[312]=25'd785;
            NN[313]=25'd5289;
            NN[314]=25'd6707;
            NN[315]=25'd10932;
            NN[316]=25'd14956;
            NN[317]=25'd14401;
            NN[318]=25'd11360;
            NN[319]=25'd7585;
            NN[320]=25'd12881;
            NN[321]=25'd12179;
            NN[322]=25'd16338;
            NN[323]=25'd10924;
            NN[324]=25'd16186;
            NN[325]=25'd19860;
            NN[326]=25'd24125;
            NN[327]=25'd29120;
            NN[328]=25'd27918;
            NN[329]=25'd19045;
            NN[330]=25'd7794;
            NN[331]=25'd3309;
            NN[332]=-25'd20;
            NN[333]=-25'd102;
            NN[334]=-25'd275;
            NN[335]=25'd0;
            NN[336]=25'd0;
            NN[337]=25'd0;
            NN[338]=25'd0;
            NN[339]=25'd0;
            NN[340]=25'd1150;
            NN[341]=25'd3041;
            NN[342]=25'd4425;
            NN[343]=25'd5297;
            NN[344]=25'd7665;
            NN[345]=25'd12034;
            NN[346]=25'd14174;
            NN[347]=25'd14291;
            NN[348]=25'd19544;
            NN[349]=25'd20034;
            NN[350]=25'd23191;
            NN[351]=25'd15455;
            NN[352]=25'd13297;
            NN[353]=25'd10017;
            NN[354]=25'd10947;
            NN[355]=25'd11330;
            NN[356]=25'd9502;
            NN[357]=25'd5758;
            NN[358]=25'd1230;
            NN[359]=25'd299;
            NN[360]=25'd23;
            NN[361]=25'd0;
            NN[362]=25'd0;
            NN[363]=25'd0;
            NN[364]=25'd0;
            NN[365]=25'd0;
            NN[366]=25'd0;
            NN[367]=25'd0;
            NN[368]=-25'd1;
            NN[369]=-25'd5;
            NN[370]=25'd52;
            NN[371]=25'd278;
            NN[372]=25'd88;
            NN[373]=25'd147;
            NN[374]=25'd384;
            NN[375]=-25'd222;
            NN[376]=25'd30;
            NN[377]=-25'd1218;
            NN[378]=25'd153;
            NN[379]=-25'd1308;
            NN[380]=-25'd1096;
            NN[381]=-25'd2025;
            NN[382]=-25'd2654;
            NN[383]=-25'd1349;
            NN[384]=25'd141;
            NN[385]=25'd574;
            NN[386]=25'd466;
            NN[387]=-25'd28;
            NN[388]=25'd0;
            NN[389]=25'd0;
            NN[390]=25'd0;
            NN[391]=25'd0;
        end
		endcase
	end
	


	
endmodule