module conv28x28(data , dPstate , core ,out);
    parameter ArraySize = 25;
    parameter   IntSize =  8;
    
    input  wire [784*IntSize-1:0] data;
    input wire [20:0] dPstate;
    input wire [ArraySize*IntSize-1:0] core;
    output wire [7:0] out;
   
    reg  [ArraySize*IntSize-1:0]  dPIn;
    
dotProduct dot1(.in1(dPIn) , .in2(core) , .out(out)); 

always @* begin
    case(dPstate)
0 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[7:0] ,data[15:8] ,data[23:16] ,0 ,0 ,data[231:224] ,data[239:232] ,data[247:240] ,0 ,0 ,data[455:448] ,data[463:456] ,data[471:464] };
end
1 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[7:0] ,data[15:8] ,data[23:16] ,data[31:24] ,0 ,data[231:224] ,data[239:232] ,data[247:240] ,data[255:248] ,0 ,data[455:448] ,data[463:456] ,data[471:464] ,data[479:472] };
end
2 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[7:0] ,data[15:8] ,data[23:16] ,data[31:24] ,data[39:32] ,data[231:224] ,data[239:232] ,data[247:240] ,data[255:248] ,data[263:256] ,data[455:448] ,data[463:456] ,data[471:464] ,data[479:472] ,data[487:480] };
end
3 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[15:8] ,data[23:16] ,data[31:24] ,data[39:32] ,data[47:40] ,data[239:232] ,data[247:240] ,data[255:248] ,data[263:256] ,data[271:264] ,data[463:456] ,data[471:464] ,data[479:472] ,data[487:480] ,data[495:488] };
end
4 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[23:16] ,data[31:24] ,data[39:32] ,data[47:40] ,data[55:48] ,data[247:240] ,data[255:248] ,data[263:256] ,data[271:264] ,data[279:272] ,data[471:464] ,data[479:472] ,data[487:480] ,data[495:488] ,data[503:496] };
end
5 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[31:24] ,data[39:32] ,data[47:40] ,data[55:48] ,data[63:56] ,data[255:248] ,data[263:256] ,data[271:264] ,data[279:272] ,data[287:280] ,data[479:472] ,data[487:480] ,data[495:488] ,data[503:496] ,data[511:504] };
end
6 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[39:32] ,data[47:40] ,data[55:48] ,data[63:56] ,data[71:64] ,data[263:256] ,data[271:264] ,data[279:272] ,data[287:280] ,data[295:288] ,data[487:480] ,data[495:488] ,data[503:496] ,data[511:504] ,data[519:512] };
end
7 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[47:40] ,data[55:48] ,data[63:56] ,data[71:64] ,data[79:72] ,data[271:264] ,data[279:272] ,data[287:280] ,data[295:288] ,data[303:296] ,data[495:488] ,data[503:496] ,data[511:504] ,data[519:512] ,data[527:520] };
end
8 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[55:48] ,data[63:56] ,data[71:64] ,data[79:72] ,data[87:80] ,data[279:272] ,data[287:280] ,data[295:288] ,data[303:296] ,data[311:304] ,data[503:496] ,data[511:504] ,data[519:512] ,data[527:520] ,data[535:528] };
end
9 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[63:56] ,data[71:64] ,data[79:72] ,data[87:80] ,data[95:88] ,data[287:280] ,data[295:288] ,data[303:296] ,data[311:304] ,data[319:312] ,data[511:504] ,data[519:512] ,data[527:520] ,data[535:528] ,data[543:536] };
end
10 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[71:64] ,data[79:72] ,data[87:80] ,data[95:88] ,data[103:96] ,data[295:288] ,data[303:296] ,data[311:304] ,data[319:312] ,data[327:320] ,data[519:512] ,data[527:520] ,data[535:528] ,data[543:536] ,data[551:544] };
end
11 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[79:72] ,data[87:80] ,data[95:88] ,data[103:96] ,data[111:104] ,data[303:296] ,data[311:304] ,data[319:312] ,data[327:320] ,data[335:328] ,data[527:520] ,data[535:528] ,data[543:536] ,data[551:544] ,data[559:552] };
end
12 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[87:80] ,data[95:88] ,data[103:96] ,data[111:104] ,data[119:112] ,data[311:304] ,data[319:312] ,data[327:320] ,data[335:328] ,data[343:336] ,data[535:528] ,data[543:536] ,data[551:544] ,data[559:552] ,data[567:560] };
end
13 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[95:88] ,data[103:96] ,data[111:104] ,data[119:112] ,data[127:120] ,data[319:312] ,data[327:320] ,data[335:328] ,data[343:336] ,data[351:344] ,data[543:536] ,data[551:544] ,data[559:552] ,data[567:560] ,data[575:568] };
end
14 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[103:96] ,data[111:104] ,data[119:112] ,data[127:120] ,data[135:128] ,data[327:320] ,data[335:328] ,data[343:336] ,data[351:344] ,data[359:352] ,data[551:544] ,data[559:552] ,data[567:560] ,data[575:568] ,data[583:576] };
end
15 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[111:104] ,data[119:112] ,data[127:120] ,data[135:128] ,data[143:136] ,data[335:328] ,data[343:336] ,data[351:344] ,data[359:352] ,data[367:360] ,data[559:552] ,data[567:560] ,data[575:568] ,data[583:576] ,data[591:584] };
end
16 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[119:112] ,data[127:120] ,data[135:128] ,data[143:136] ,data[151:144] ,data[343:336] ,data[351:344] ,data[359:352] ,data[367:360] ,data[375:368] ,data[567:560] ,data[575:568] ,data[583:576] ,data[591:584] ,data[599:592] };
end
17 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[127:120] ,data[135:128] ,data[143:136] ,data[151:144] ,data[159:152] ,data[351:344] ,data[359:352] ,data[367:360] ,data[375:368] ,data[383:376] ,data[575:568] ,data[583:576] ,data[591:584] ,data[599:592] ,data[607:600] };
end
18 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[135:128] ,data[143:136] ,data[151:144] ,data[159:152] ,data[167:160] ,data[359:352] ,data[367:360] ,data[375:368] ,data[383:376] ,data[391:384] ,data[583:576] ,data[591:584] ,data[599:592] ,data[607:600] ,data[615:608] };
end
19 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[143:136] ,data[151:144] ,data[159:152] ,data[167:160] ,data[175:168] ,data[367:360] ,data[375:368] ,data[383:376] ,data[391:384] ,data[399:392] ,data[591:584] ,data[599:592] ,data[607:600] ,data[615:608] ,data[623:616] };
end
20 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[151:144] ,data[159:152] ,data[167:160] ,data[175:168] ,data[183:176] ,data[375:368] ,data[383:376] ,data[391:384] ,data[399:392] ,data[407:400] ,data[599:592] ,data[607:600] ,data[615:608] ,data[623:616] ,data[631:624] };
end
21 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[159:152] ,data[167:160] ,data[175:168] ,data[183:176] ,data[191:184] ,data[383:376] ,data[391:384] ,data[399:392] ,data[407:400] ,data[415:408] ,data[607:600] ,data[615:608] ,data[623:616] ,data[631:624] ,data[639:632] };
end
22 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[167:160] ,data[175:168] ,data[183:176] ,data[191:184] ,data[199:192] ,data[391:384] ,data[399:392] ,data[407:400] ,data[415:408] ,data[423:416] ,data[615:608] ,data[623:616] ,data[631:624] ,data[639:632] ,data[647:640] };
end
23 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[175:168] ,data[183:176] ,data[191:184] ,data[199:192] ,data[207:200] ,data[399:392] ,data[407:400] ,data[415:408] ,data[423:416] ,data[431:424] ,data[623:616] ,data[631:624] ,data[639:632] ,data[647:640] ,data[655:648] };
end
24 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[183:176] ,data[191:184] ,data[199:192] ,data[207:200] ,data[215:208] ,data[407:400] ,data[415:408] ,data[423:416] ,data[431:424] ,data[439:432] ,data[631:624] ,data[639:632] ,data[647:640] ,data[655:648] ,data[663:656] };
end
25 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[191:184] ,data[199:192] ,data[207:200] ,data[215:208] ,data[223:216] ,data[415:408] ,data[423:416] ,data[431:424] ,data[439:432] ,data[447:440] ,data[639:632] ,data[647:640] ,data[655:648] ,data[663:656] ,data[671:664] };
end
26 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[199:192] ,data[207:200] ,data[215:208] ,data[223:216] ,0 ,data[423:416] ,data[431:424] ,data[439:432] ,data[447:440] ,0 ,data[647:640] ,data[655:648] ,data[663:656] ,data[671:664] ,0 };
end
27 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[207:200] ,data[215:208] ,data[223:216] ,0 ,0 ,data[431:424] ,data[439:432] ,data[447:440] ,0 ,0 ,data[655:648] ,data[663:656] ,data[671:664] ,0 ,0 };
end
28 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,0 ,data[7:0] ,data[15:8] ,data[23:16] ,0 ,0 ,data[231:224] ,data[239:232] ,data[247:240] ,0 ,0 ,data[455:448] ,data[463:456] ,data[471:464] ,0 ,0 ,data[679:672] ,data[687:680] ,data[695:688] };
end
29 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,0 ,data[7:0] ,data[15:8] ,data[23:16] ,data[31:24] ,0 ,data[231:224] ,data[239:232] ,data[247:240] ,data[255:248] ,0 ,data[455:448] ,data[463:456] ,data[471:464] ,data[479:472] ,0 ,data[679:672] ,data[687:680] ,data[695:688] ,data[703:696] };
end
30 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[7:0] ,data[15:8] ,data[23:16] ,data[31:24] ,data[39:32] ,data[231:224] ,data[239:232] ,data[247:240] ,data[255:248] ,data[263:256] ,data[455:448] ,data[463:456] ,data[471:464] ,data[479:472] ,data[487:480] ,data[679:672] ,data[687:680] ,data[695:688] ,data[703:696] ,data[711:704] };
end
31 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[15:8] ,data[23:16] ,data[31:24] ,data[39:32] ,data[47:40] ,data[239:232] ,data[247:240] ,data[255:248] ,data[263:256] ,data[271:264] ,data[463:456] ,data[471:464] ,data[479:472] ,data[487:480] ,data[495:488] ,data[687:680] ,data[695:688] ,data[703:696] ,data[711:704] ,data[719:712] };
end
32 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[23:16] ,data[31:24] ,data[39:32] ,data[47:40] ,data[55:48] ,data[247:240] ,data[255:248] ,data[263:256] ,data[271:264] ,data[279:272] ,data[471:464] ,data[479:472] ,data[487:480] ,data[495:488] ,data[503:496] ,data[695:688] ,data[703:696] ,data[711:704] ,data[719:712] ,data[727:720] };
end
33 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[31:24] ,data[39:32] ,data[47:40] ,data[55:48] ,data[63:56] ,data[255:248] ,data[263:256] ,data[271:264] ,data[279:272] ,data[287:280] ,data[479:472] ,data[487:480] ,data[495:488] ,data[503:496] ,data[511:504] ,data[703:696] ,data[711:704] ,data[719:712] ,data[727:720] ,data[735:728] };
end
34 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[39:32] ,data[47:40] ,data[55:48] ,data[63:56] ,data[71:64] ,data[263:256] ,data[271:264] ,data[279:272] ,data[287:280] ,data[295:288] ,data[487:480] ,data[495:488] ,data[503:496] ,data[511:504] ,data[519:512] ,data[711:704] ,data[719:712] ,data[727:720] ,data[735:728] ,data[743:736] };
end
35 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[47:40] ,data[55:48] ,data[63:56] ,data[71:64] ,data[79:72] ,data[271:264] ,data[279:272] ,data[287:280] ,data[295:288] ,data[303:296] ,data[495:488] ,data[503:496] ,data[511:504] ,data[519:512] ,data[527:520] ,data[719:712] ,data[727:720] ,data[735:728] ,data[743:736] ,data[751:744] };
end
36 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[55:48] ,data[63:56] ,data[71:64] ,data[79:72] ,data[87:80] ,data[279:272] ,data[287:280] ,data[295:288] ,data[303:296] ,data[311:304] ,data[503:496] ,data[511:504] ,data[519:512] ,data[527:520] ,data[535:528] ,data[727:720] ,data[735:728] ,data[743:736] ,data[751:744] ,data[759:752] };
end
37 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[63:56] ,data[71:64] ,data[79:72] ,data[87:80] ,data[95:88] ,data[287:280] ,data[295:288] ,data[303:296] ,data[311:304] ,data[319:312] ,data[511:504] ,data[519:512] ,data[527:520] ,data[535:528] ,data[543:536] ,data[735:728] ,data[743:736] ,data[751:744] ,data[759:752] ,data[767:760] };
end
38 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[71:64] ,data[79:72] ,data[87:80] ,data[95:88] ,data[103:96] ,data[295:288] ,data[303:296] ,data[311:304] ,data[319:312] ,data[327:320] ,data[519:512] ,data[527:520] ,data[535:528] ,data[543:536] ,data[551:544] ,data[743:736] ,data[751:744] ,data[759:752] ,data[767:760] ,data[775:768] };
end
39 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[79:72] ,data[87:80] ,data[95:88] ,data[103:96] ,data[111:104] ,data[303:296] ,data[311:304] ,data[319:312] ,data[327:320] ,data[335:328] ,data[527:520] ,data[535:528] ,data[543:536] ,data[551:544] ,data[559:552] ,data[751:744] ,data[759:752] ,data[767:760] ,data[775:768] ,data[783:776] };
end
40 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[87:80] ,data[95:88] ,data[103:96] ,data[111:104] ,data[119:112] ,data[311:304] ,data[319:312] ,data[327:320] ,data[335:328] ,data[343:336] ,data[535:528] ,data[543:536] ,data[551:544] ,data[559:552] ,data[567:560] ,data[759:752] ,data[767:760] ,data[775:768] ,data[783:776] ,data[791:784] };
end
41 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[95:88] ,data[103:96] ,data[111:104] ,data[119:112] ,data[127:120] ,data[319:312] ,data[327:320] ,data[335:328] ,data[343:336] ,data[351:344] ,data[543:536] ,data[551:544] ,data[559:552] ,data[567:560] ,data[575:568] ,data[767:760] ,data[775:768] ,data[783:776] ,data[791:784] ,data[799:792] };
end
42 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[103:96] ,data[111:104] ,data[119:112] ,data[127:120] ,data[135:128] ,data[327:320] ,data[335:328] ,data[343:336] ,data[351:344] ,data[359:352] ,data[551:544] ,data[559:552] ,data[567:560] ,data[575:568] ,data[583:576] ,data[775:768] ,data[783:776] ,data[791:784] ,data[799:792] ,data[807:800] };
end
43 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[111:104] ,data[119:112] ,data[127:120] ,data[135:128] ,data[143:136] ,data[335:328] ,data[343:336] ,data[351:344] ,data[359:352] ,data[367:360] ,data[559:552] ,data[567:560] ,data[575:568] ,data[583:576] ,data[591:584] ,data[783:776] ,data[791:784] ,data[799:792] ,data[807:800] ,data[815:808] };
end
44 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[119:112] ,data[127:120] ,data[135:128] ,data[143:136] ,data[151:144] ,data[343:336] ,data[351:344] ,data[359:352] ,data[367:360] ,data[375:368] ,data[567:560] ,data[575:568] ,data[583:576] ,data[591:584] ,data[599:592] ,data[791:784] ,data[799:792] ,data[807:800] ,data[815:808] ,data[823:816] };
end
45 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[127:120] ,data[135:128] ,data[143:136] ,data[151:144] ,data[159:152] ,data[351:344] ,data[359:352] ,data[367:360] ,data[375:368] ,data[383:376] ,data[575:568] ,data[583:576] ,data[591:584] ,data[599:592] ,data[607:600] ,data[799:792] ,data[807:800] ,data[815:808] ,data[823:816] ,data[831:824] };
end
46 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[135:128] ,data[143:136] ,data[151:144] ,data[159:152] ,data[167:160] ,data[359:352] ,data[367:360] ,data[375:368] ,data[383:376] ,data[391:384] ,data[583:576] ,data[591:584] ,data[599:592] ,data[607:600] ,data[615:608] ,data[807:800] ,data[815:808] ,data[823:816] ,data[831:824] ,data[839:832] };
end
47 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[143:136] ,data[151:144] ,data[159:152] ,data[167:160] ,data[175:168] ,data[367:360] ,data[375:368] ,data[383:376] ,data[391:384] ,data[399:392] ,data[591:584] ,data[599:592] ,data[607:600] ,data[615:608] ,data[623:616] ,data[815:808] ,data[823:816] ,data[831:824] ,data[839:832] ,data[847:840] };
end
48 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[151:144] ,data[159:152] ,data[167:160] ,data[175:168] ,data[183:176] ,data[375:368] ,data[383:376] ,data[391:384] ,data[399:392] ,data[407:400] ,data[599:592] ,data[607:600] ,data[615:608] ,data[623:616] ,data[631:624] ,data[823:816] ,data[831:824] ,data[839:832] ,data[847:840] ,data[855:848] };
end
49 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[159:152] ,data[167:160] ,data[175:168] ,data[183:176] ,data[191:184] ,data[383:376] ,data[391:384] ,data[399:392] ,data[407:400] ,data[415:408] ,data[607:600] ,data[615:608] ,data[623:616] ,data[631:624] ,data[639:632] ,data[831:824] ,data[839:832] ,data[847:840] ,data[855:848] ,data[863:856] };
end
50 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[167:160] ,data[175:168] ,data[183:176] ,data[191:184] ,data[199:192] ,data[391:384] ,data[399:392] ,data[407:400] ,data[415:408] ,data[423:416] ,data[615:608] ,data[623:616] ,data[631:624] ,data[639:632] ,data[647:640] ,data[839:832] ,data[847:840] ,data[855:848] ,data[863:856] ,data[871:864] };
end
51 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[175:168] ,data[183:176] ,data[191:184] ,data[199:192] ,data[207:200] ,data[399:392] ,data[407:400] ,data[415:408] ,data[423:416] ,data[431:424] ,data[623:616] ,data[631:624] ,data[639:632] ,data[647:640] ,data[655:648] ,data[847:840] ,data[855:848] ,data[863:856] ,data[871:864] ,data[879:872] };
end
52 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[183:176] ,data[191:184] ,data[199:192] ,data[207:200] ,data[215:208] ,data[407:400] ,data[415:408] ,data[423:416] ,data[431:424] ,data[439:432] ,data[631:624] ,data[639:632] ,data[647:640] ,data[655:648] ,data[663:656] ,data[855:848] ,data[863:856] ,data[871:864] ,data[879:872] ,data[887:880] };
end
53 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[191:184] ,data[199:192] ,data[207:200] ,data[215:208] ,data[223:216] ,data[415:408] ,data[423:416] ,data[431:424] ,data[439:432] ,data[447:440] ,data[639:632] ,data[647:640] ,data[655:648] ,data[663:656] ,data[671:664] ,data[863:856] ,data[871:864] ,data[879:872] ,data[887:880] ,data[895:888] };
end
54 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[199:192] ,data[207:200] ,data[215:208] ,data[223:216] ,0 ,data[423:416] ,data[431:424] ,data[439:432] ,data[447:440] ,0 ,data[647:640] ,data[655:648] ,data[663:656] ,data[671:664] ,0 ,data[871:864] ,data[879:872] ,data[887:880] ,data[895:888] ,0 };
end
55 :begin
 dPIn = {0 ,0 ,0 ,0 ,0 ,data[207:200] ,data[215:208] ,data[223:216] ,0 ,0 ,data[431:424] ,data[439:432] ,data[447:440] ,0 ,0 ,data[655:648] ,data[663:656] ,data[671:664] ,0 ,0 ,data[879:872] ,data[887:880] ,data[895:888] ,0 ,0 };
end
56 :begin
 dPIn = {0 ,0 ,data[7:0] ,data[15:8] ,data[23:16] ,0 ,0 ,data[231:224] ,data[239:232] ,data[247:240] ,0 ,0 ,data[455:448] ,data[463:456] ,data[471:464] ,0 ,0 ,data[679:672] ,data[687:680] ,data[695:688] ,0 ,0 ,data[903:896] ,data[911:904] ,data[919:912] };
end
57 :begin
 dPIn = {0 ,data[7:0] ,data[15:8] ,data[23:16] ,data[31:24] ,0 ,data[231:224] ,data[239:232] ,data[247:240] ,data[255:248] ,0 ,data[455:448] ,data[463:456] ,data[471:464] ,data[479:472] ,0 ,data[679:672] ,data[687:680] ,data[695:688] ,data[703:696] ,0 ,data[903:896] ,data[911:904] ,data[919:912] ,data[927:920] };
end
58 :begin
 dPIn = {data[7:0] ,data[15:8] ,data[23:16] ,data[31:24] ,data[39:32] ,data[231:224] ,data[239:232] ,data[247:240] ,data[255:248] ,data[263:256] ,data[455:448] ,data[463:456] ,data[471:464] ,data[479:472] ,data[487:480] ,data[679:672] ,data[687:680] ,data[695:688] ,data[703:696] ,data[711:704] ,data[903:896] ,data[911:904] ,data[919:912] ,data[927:920] ,data[935:928] };
end
59 :begin
 dPIn = {data[15:8] ,data[23:16] ,data[31:24] ,data[39:32] ,data[47:40] ,data[239:232] ,data[247:240] ,data[255:248] ,data[263:256] ,data[271:264] ,data[463:456] ,data[471:464] ,data[479:472] ,data[487:480] ,data[495:488] ,data[687:680] ,data[695:688] ,data[703:696] ,data[711:704] ,data[719:712] ,data[911:904] ,data[919:912] ,data[927:920] ,data[935:928] ,data[943:936] };
end
60 :begin
 dPIn = {data[23:16] ,data[31:24] ,data[39:32] ,data[47:40] ,data[55:48] ,data[247:240] ,data[255:248] ,data[263:256] ,data[271:264] ,data[279:272] ,data[471:464] ,data[479:472] ,data[487:480] ,data[495:488] ,data[503:496] ,data[695:688] ,data[703:696] ,data[711:704] ,data[719:712] ,data[727:720] ,data[919:912] ,data[927:920] ,data[935:928] ,data[943:936] ,data[951:944] };
end
61 :begin
 dPIn = {data[31:24] ,data[39:32] ,data[47:40] ,data[55:48] ,data[63:56] ,data[255:248] ,data[263:256] ,data[271:264] ,data[279:272] ,data[287:280] ,data[479:472] ,data[487:480] ,data[495:488] ,data[503:496] ,data[511:504] ,data[703:696] ,data[711:704] ,data[719:712] ,data[727:720] ,data[735:728] ,data[927:920] ,data[935:928] ,data[943:936] ,data[951:944] ,data[959:952] };
end
62 :begin
 dPIn = {data[39:32] ,data[47:40] ,data[55:48] ,data[63:56] ,data[71:64] ,data[263:256] ,data[271:264] ,data[279:272] ,data[287:280] ,data[295:288] ,data[487:480] ,data[495:488] ,data[503:496] ,data[511:504] ,data[519:512] ,data[711:704] ,data[719:712] ,data[727:720] ,data[735:728] ,data[743:736] ,data[935:928] ,data[943:936] ,data[951:944] ,data[959:952] ,data[967:960] };
end
63 :begin
 dPIn = {data[47:40] ,data[55:48] ,data[63:56] ,data[71:64] ,data[79:72] ,data[271:264] ,data[279:272] ,data[287:280] ,data[295:288] ,data[303:296] ,data[495:488] ,data[503:496] ,data[511:504] ,data[519:512] ,data[527:520] ,data[719:712] ,data[727:720] ,data[735:728] ,data[743:736] ,data[751:744] ,data[943:936] ,data[951:944] ,data[959:952] ,data[967:960] ,data[975:968] };
end
64 :begin
 dPIn = {data[55:48] ,data[63:56] ,data[71:64] ,data[79:72] ,data[87:80] ,data[279:272] ,data[287:280] ,data[295:288] ,data[303:296] ,data[311:304] ,data[503:496] ,data[511:504] ,data[519:512] ,data[527:520] ,data[535:528] ,data[727:720] ,data[735:728] ,data[743:736] ,data[751:744] ,data[759:752] ,data[951:944] ,data[959:952] ,data[967:960] ,data[975:968] ,data[983:976] };
end
65 :begin
 dPIn = {data[63:56] ,data[71:64] ,data[79:72] ,data[87:80] ,data[95:88] ,data[287:280] ,data[295:288] ,data[303:296] ,data[311:304] ,data[319:312] ,data[511:504] ,data[519:512] ,data[527:520] ,data[535:528] ,data[543:536] ,data[735:728] ,data[743:736] ,data[751:744] ,data[759:752] ,data[767:760] ,data[959:952] ,data[967:960] ,data[975:968] ,data[983:976] ,data[991:984] };
end
66 :begin
 dPIn = {data[71:64] ,data[79:72] ,data[87:80] ,data[95:88] ,data[103:96] ,data[295:288] ,data[303:296] ,data[311:304] ,data[319:312] ,data[327:320] ,data[519:512] ,data[527:520] ,data[535:528] ,data[543:536] ,data[551:544] ,data[743:736] ,data[751:744] ,data[759:752] ,data[767:760] ,data[775:768] ,data[967:960] ,data[975:968] ,data[983:976] ,data[991:984] ,data[999:992] };
end
67 :begin
 dPIn = {data[79:72] ,data[87:80] ,data[95:88] ,data[103:96] ,data[111:104] ,data[303:296] ,data[311:304] ,data[319:312] ,data[327:320] ,data[335:328] ,data[527:520] ,data[535:528] ,data[543:536] ,data[551:544] ,data[559:552] ,data[751:744] ,data[759:752] ,data[767:760] ,data[775:768] ,data[783:776] ,data[975:968] ,data[983:976] ,data[991:984] ,data[999:992] ,data[1007:1000] };
end
68 :begin
 dPIn = {data[87:80] ,data[95:88] ,data[103:96] ,data[111:104] ,data[119:112] ,data[311:304] ,data[319:312] ,data[327:320] ,data[335:328] ,data[343:336] ,data[535:528] ,data[543:536] ,data[551:544] ,data[559:552] ,data[567:560] ,data[759:752] ,data[767:760] ,data[775:768] ,data[783:776] ,data[791:784] ,data[983:976] ,data[991:984] ,data[999:992] ,data[1007:1000] ,data[1015:1008] };
end
69 :begin
 dPIn = {data[95:88] ,data[103:96] ,data[111:104] ,data[119:112] ,data[127:120] ,data[319:312] ,data[327:320] ,data[335:328] ,data[343:336] ,data[351:344] ,data[543:536] ,data[551:544] ,data[559:552] ,data[567:560] ,data[575:568] ,data[767:760] ,data[775:768] ,data[783:776] ,data[791:784] ,data[799:792] ,data[991:984] ,data[999:992] ,data[1007:1000] ,data[1015:1008] ,data[1023:1016] };
end
70 :begin
 dPIn = {data[103:96] ,data[111:104] ,data[119:112] ,data[127:120] ,data[135:128] ,data[327:320] ,data[335:328] ,data[343:336] ,data[351:344] ,data[359:352] ,data[551:544] ,data[559:552] ,data[567:560] ,data[575:568] ,data[583:576] ,data[775:768] ,data[783:776] ,data[791:784] ,data[799:792] ,data[807:800] ,data[999:992] ,data[1007:1000] ,data[1015:1008] ,data[1023:1016] ,data[1031:1024] };
end
71 :begin
 dPIn = {data[111:104] ,data[119:112] ,data[127:120] ,data[135:128] ,data[143:136] ,data[335:328] ,data[343:336] ,data[351:344] ,data[359:352] ,data[367:360] ,data[559:552] ,data[567:560] ,data[575:568] ,data[583:576] ,data[591:584] ,data[783:776] ,data[791:784] ,data[799:792] ,data[807:800] ,data[815:808] ,data[1007:1000] ,data[1015:1008] ,data[1023:1016] ,data[1031:1024] ,data[1039:1032] };
end
72 :begin
 dPIn = {data[119:112] ,data[127:120] ,data[135:128] ,data[143:136] ,data[151:144] ,data[343:336] ,data[351:344] ,data[359:352] ,data[367:360] ,data[375:368] ,data[567:560] ,data[575:568] ,data[583:576] ,data[591:584] ,data[599:592] ,data[791:784] ,data[799:792] ,data[807:800] ,data[815:808] ,data[823:816] ,data[1015:1008] ,data[1023:1016] ,data[1031:1024] ,data[1039:1032] ,data[1047:1040] };
end
73 :begin
 dPIn = {data[127:120] ,data[135:128] ,data[143:136] ,data[151:144] ,data[159:152] ,data[351:344] ,data[359:352] ,data[367:360] ,data[375:368] ,data[383:376] ,data[575:568] ,data[583:576] ,data[591:584] ,data[599:592] ,data[607:600] ,data[799:792] ,data[807:800] ,data[815:808] ,data[823:816] ,data[831:824] ,data[1023:1016] ,data[1031:1024] ,data[1039:1032] ,data[1047:1040] ,data[1055:1048] };
end
74 :begin
 dPIn = {data[135:128] ,data[143:136] ,data[151:144] ,data[159:152] ,data[167:160] ,data[359:352] ,data[367:360] ,data[375:368] ,data[383:376] ,data[391:384] ,data[583:576] ,data[591:584] ,data[599:592] ,data[607:600] ,data[615:608] ,data[807:800] ,data[815:808] ,data[823:816] ,data[831:824] ,data[839:832] ,data[1031:1024] ,data[1039:1032] ,data[1047:1040] ,data[1055:1048] ,data[1063:1056] };
end
75 :begin
 dPIn = {data[143:136] ,data[151:144] ,data[159:152] ,data[167:160] ,data[175:168] ,data[367:360] ,data[375:368] ,data[383:376] ,data[391:384] ,data[399:392] ,data[591:584] ,data[599:592] ,data[607:600] ,data[615:608] ,data[623:616] ,data[815:808] ,data[823:816] ,data[831:824] ,data[839:832] ,data[847:840] ,data[1039:1032] ,data[1047:1040] ,data[1055:1048] ,data[1063:1056] ,data[1071:1064] };
end
76 :begin
 dPIn = {data[151:144] ,data[159:152] ,data[167:160] ,data[175:168] ,data[183:176] ,data[375:368] ,data[383:376] ,data[391:384] ,data[399:392] ,data[407:400] ,data[599:592] ,data[607:600] ,data[615:608] ,data[623:616] ,data[631:624] ,data[823:816] ,data[831:824] ,data[839:832] ,data[847:840] ,data[855:848] ,data[1047:1040] ,data[1055:1048] ,data[1063:1056] ,data[1071:1064] ,data[1079:1072] };
end
77 :begin
 dPIn = {data[159:152] ,data[167:160] ,data[175:168] ,data[183:176] ,data[191:184] ,data[383:376] ,data[391:384] ,data[399:392] ,data[407:400] ,data[415:408] ,data[607:600] ,data[615:608] ,data[623:616] ,data[631:624] ,data[639:632] ,data[831:824] ,data[839:832] ,data[847:840] ,data[855:848] ,data[863:856] ,data[1055:1048] ,data[1063:1056] ,data[1071:1064] ,data[1079:1072] ,data[1087:1080] };
end
78 :begin
 dPIn = {data[167:160] ,data[175:168] ,data[183:176] ,data[191:184] ,data[199:192] ,data[391:384] ,data[399:392] ,data[407:400] ,data[415:408] ,data[423:416] ,data[615:608] ,data[623:616] ,data[631:624] ,data[639:632] ,data[647:640] ,data[839:832] ,data[847:840] ,data[855:848] ,data[863:856] ,data[871:864] ,data[1063:1056] ,data[1071:1064] ,data[1079:1072] ,data[1087:1080] ,data[1095:1088] };
end
79 :begin
 dPIn = {data[175:168] ,data[183:176] ,data[191:184] ,data[199:192] ,data[207:200] ,data[399:392] ,data[407:400] ,data[415:408] ,data[423:416] ,data[431:424] ,data[623:616] ,data[631:624] ,data[639:632] ,data[647:640] ,data[655:648] ,data[847:840] ,data[855:848] ,data[863:856] ,data[871:864] ,data[879:872] ,data[1071:1064] ,data[1079:1072] ,data[1087:1080] ,data[1095:1088] ,data[1103:1096] };
end
80 :begin
 dPIn = {data[183:176] ,data[191:184] ,data[199:192] ,data[207:200] ,data[215:208] ,data[407:400] ,data[415:408] ,data[423:416] ,data[431:424] ,data[439:432] ,data[631:624] ,data[639:632] ,data[647:640] ,data[655:648] ,data[663:656] ,data[855:848] ,data[863:856] ,data[871:864] ,data[879:872] ,data[887:880] ,data[1079:1072] ,data[1087:1080] ,data[1095:1088] ,data[1103:1096] ,data[1111:1104] };
end
81 :begin
 dPIn = {data[191:184] ,data[199:192] ,data[207:200] ,data[215:208] ,data[223:216] ,data[415:408] ,data[423:416] ,data[431:424] ,data[439:432] ,data[447:440] ,data[639:632] ,data[647:640] ,data[655:648] ,data[663:656] ,data[671:664] ,data[863:856] ,data[871:864] ,data[879:872] ,data[887:880] ,data[895:888] ,data[1087:1080] ,data[1095:1088] ,data[1103:1096] ,data[1111:1104] ,data[1119:1112] };
end
82 :begin
 dPIn = {data[199:192] ,data[207:200] ,data[215:208] ,data[223:216] ,0 ,data[423:416] ,data[431:424] ,data[439:432] ,data[447:440] ,0 ,data[647:640] ,data[655:648] ,data[663:656] ,data[671:664] ,0 ,data[871:864] ,data[879:872] ,data[887:880] ,data[895:888] ,0 ,data[1095:1088] ,data[1103:1096] ,data[1111:1104] ,data[1119:1112] ,0 };
end
83 :begin
 dPIn = {data[207:200] ,data[215:208] ,data[223:216] ,0 ,0 ,data[431:424] ,data[439:432] ,data[447:440] ,0 ,0 ,data[655:648] ,data[663:656] ,data[671:664] ,0 ,0 ,data[879:872] ,data[887:880] ,data[895:888] ,0 ,0 ,data[1103:1096] ,data[1111:1104] ,data[1119:1112] ,0 ,0 };
end
84 :begin
 dPIn = {0 ,0 ,data[231:224] ,data[239:232] ,data[247:240] ,0 ,0 ,data[455:448] ,data[463:456] ,data[471:464] ,0 ,0 ,data[679:672] ,data[687:680] ,data[695:688] ,0 ,0 ,data[903:896] ,data[911:904] ,data[919:912] ,0 ,0 ,data[1127:1120] ,data[1135:1128] ,data[1143:1136] };
end
85 :begin
 dPIn = {0 ,data[231:224] ,data[239:232] ,data[247:240] ,data[255:248] ,0 ,data[455:448] ,data[463:456] ,data[471:464] ,data[479:472] ,0 ,data[679:672] ,data[687:680] ,data[695:688] ,data[703:696] ,0 ,data[903:896] ,data[911:904] ,data[919:912] ,data[927:920] ,0 ,data[1127:1120] ,data[1135:1128] ,data[1143:1136] ,data[1151:1144] };
end
86 :begin
 dPIn = {data[231:224] ,data[239:232] ,data[247:240] ,data[255:248] ,data[263:256] ,data[455:448] ,data[463:456] ,data[471:464] ,data[479:472] ,data[487:480] ,data[679:672] ,data[687:680] ,data[695:688] ,data[703:696] ,data[711:704] ,data[903:896] ,data[911:904] ,data[919:912] ,data[927:920] ,data[935:928] ,data[1127:1120] ,data[1135:1128] ,data[1143:1136] ,data[1151:1144] ,data[1159:1152] };
end
87 :begin
 dPIn = {data[239:232] ,data[247:240] ,data[255:248] ,data[263:256] ,data[271:264] ,data[463:456] ,data[471:464] ,data[479:472] ,data[487:480] ,data[495:488] ,data[687:680] ,data[695:688] ,data[703:696] ,data[711:704] ,data[719:712] ,data[911:904] ,data[919:912] ,data[927:920] ,data[935:928] ,data[943:936] ,data[1135:1128] ,data[1143:1136] ,data[1151:1144] ,data[1159:1152] ,data[1167:1160] };
end
88 :begin
 dPIn = {data[247:240] ,data[255:248] ,data[263:256] ,data[271:264] ,data[279:272] ,data[471:464] ,data[479:472] ,data[487:480] ,data[495:488] ,data[503:496] ,data[695:688] ,data[703:696] ,data[711:704] ,data[719:712] ,data[727:720] ,data[919:912] ,data[927:920] ,data[935:928] ,data[943:936] ,data[951:944] ,data[1143:1136] ,data[1151:1144] ,data[1159:1152] ,data[1167:1160] ,data[1175:1168] };
end
89 :begin
 dPIn = {data[255:248] ,data[263:256] ,data[271:264] ,data[279:272] ,data[287:280] ,data[479:472] ,data[487:480] ,data[495:488] ,data[503:496] ,data[511:504] ,data[703:696] ,data[711:704] ,data[719:712] ,data[727:720] ,data[735:728] ,data[927:920] ,data[935:928] ,data[943:936] ,data[951:944] ,data[959:952] ,data[1151:1144] ,data[1159:1152] ,data[1167:1160] ,data[1175:1168] ,data[1183:1176] };
end
90 :begin
 dPIn = {data[263:256] ,data[271:264] ,data[279:272] ,data[287:280] ,data[295:288] ,data[487:480] ,data[495:488] ,data[503:496] ,data[511:504] ,data[519:512] ,data[711:704] ,data[719:712] ,data[727:720] ,data[735:728] ,data[743:736] ,data[935:928] ,data[943:936] ,data[951:944] ,data[959:952] ,data[967:960] ,data[1159:1152] ,data[1167:1160] ,data[1175:1168] ,data[1183:1176] ,data[1191:1184] };
end
91 :begin
 dPIn = {data[271:264] ,data[279:272] ,data[287:280] ,data[295:288] ,data[303:296] ,data[495:488] ,data[503:496] ,data[511:504] ,data[519:512] ,data[527:520] ,data[719:712] ,data[727:720] ,data[735:728] ,data[743:736] ,data[751:744] ,data[943:936] ,data[951:944] ,data[959:952] ,data[967:960] ,data[975:968] ,data[1167:1160] ,data[1175:1168] ,data[1183:1176] ,data[1191:1184] ,data[1199:1192] };
end
92 :begin
 dPIn = {data[279:272] ,data[287:280] ,data[295:288] ,data[303:296] ,data[311:304] ,data[503:496] ,data[511:504] ,data[519:512] ,data[527:520] ,data[535:528] ,data[727:720] ,data[735:728] ,data[743:736] ,data[751:744] ,data[759:752] ,data[951:944] ,data[959:952] ,data[967:960] ,data[975:968] ,data[983:976] ,data[1175:1168] ,data[1183:1176] ,data[1191:1184] ,data[1199:1192] ,data[1207:1200] };
end
93 :begin
 dPIn = {data[287:280] ,data[295:288] ,data[303:296] ,data[311:304] ,data[319:312] ,data[511:504] ,data[519:512] ,data[527:520] ,data[535:528] ,data[543:536] ,data[735:728] ,data[743:736] ,data[751:744] ,data[759:752] ,data[767:760] ,data[959:952] ,data[967:960] ,data[975:968] ,data[983:976] ,data[991:984] ,data[1183:1176] ,data[1191:1184] ,data[1199:1192] ,data[1207:1200] ,data[1215:1208] };
end
94 :begin
 dPIn = {data[295:288] ,data[303:296] ,data[311:304] ,data[319:312] ,data[327:320] ,data[519:512] ,data[527:520] ,data[535:528] ,data[543:536] ,data[551:544] ,data[743:736] ,data[751:744] ,data[759:752] ,data[767:760] ,data[775:768] ,data[967:960] ,data[975:968] ,data[983:976] ,data[991:984] ,data[999:992] ,data[1191:1184] ,data[1199:1192] ,data[1207:1200] ,data[1215:1208] ,data[1223:1216] };
end
95 :begin
 dPIn = {data[303:296] ,data[311:304] ,data[319:312] ,data[327:320] ,data[335:328] ,data[527:520] ,data[535:528] ,data[543:536] ,data[551:544] ,data[559:552] ,data[751:744] ,data[759:752] ,data[767:760] ,data[775:768] ,data[783:776] ,data[975:968] ,data[983:976] ,data[991:984] ,data[999:992] ,data[1007:1000] ,data[1199:1192] ,data[1207:1200] ,data[1215:1208] ,data[1223:1216] ,data[1231:1224] };
end
96 :begin
 dPIn = {data[311:304] ,data[319:312] ,data[327:320] ,data[335:328] ,data[343:336] ,data[535:528] ,data[543:536] ,data[551:544] ,data[559:552] ,data[567:560] ,data[759:752] ,data[767:760] ,data[775:768] ,data[783:776] ,data[791:784] ,data[983:976] ,data[991:984] ,data[999:992] ,data[1007:1000] ,data[1015:1008] ,data[1207:1200] ,data[1215:1208] ,data[1223:1216] ,data[1231:1224] ,data[1239:1232] };
end
97 :begin
 dPIn = {data[319:312] ,data[327:320] ,data[335:328] ,data[343:336] ,data[351:344] ,data[543:536] ,data[551:544] ,data[559:552] ,data[567:560] ,data[575:568] ,data[767:760] ,data[775:768] ,data[783:776] ,data[791:784] ,data[799:792] ,data[991:984] ,data[999:992] ,data[1007:1000] ,data[1015:1008] ,data[1023:1016] ,data[1215:1208] ,data[1223:1216] ,data[1231:1224] ,data[1239:1232] ,data[1247:1240] };
end
98 :begin
 dPIn = {data[327:320] ,data[335:328] ,data[343:336] ,data[351:344] ,data[359:352] ,data[551:544] ,data[559:552] ,data[567:560] ,data[575:568] ,data[583:576] ,data[775:768] ,data[783:776] ,data[791:784] ,data[799:792] ,data[807:800] ,data[999:992] ,data[1007:1000] ,data[1015:1008] ,data[1023:1016] ,data[1031:1024] ,data[1223:1216] ,data[1231:1224] ,data[1239:1232] ,data[1247:1240] ,data[1255:1248] };
end
99 :begin
 dPIn = {data[335:328] ,data[343:336] ,data[351:344] ,data[359:352] ,data[367:360] ,data[559:552] ,data[567:560] ,data[575:568] ,data[583:576] ,data[591:584] ,data[783:776] ,data[791:784] ,data[799:792] ,data[807:800] ,data[815:808] ,data[1007:1000] ,data[1015:1008] ,data[1023:1016] ,data[1031:1024] ,data[1039:1032] ,data[1231:1224] ,data[1239:1232] ,data[1247:1240] ,data[1255:1248] ,data[1263:1256] };
end
100 :begin
 dPIn = {data[343:336] ,data[351:344] ,data[359:352] ,data[367:360] ,data[375:368] ,data[567:560] ,data[575:568] ,data[583:576] ,data[591:584] ,data[599:592] ,data[791:784] ,data[799:792] ,data[807:800] ,data[815:808] ,data[823:816] ,data[1015:1008] ,data[1023:1016] ,data[1031:1024] ,data[1039:1032] ,data[1047:1040] ,data[1239:1232] ,data[1247:1240] ,data[1255:1248] ,data[1263:1256] ,data[1271:1264] };
end
101 :begin
 dPIn = {data[351:344] ,data[359:352] ,data[367:360] ,data[375:368] ,data[383:376] ,data[575:568] ,data[583:576] ,data[591:584] ,data[599:592] ,data[607:600] ,data[799:792] ,data[807:800] ,data[815:808] ,data[823:816] ,data[831:824] ,data[1023:1016] ,data[1031:1024] ,data[1039:1032] ,data[1047:1040] ,data[1055:1048] ,data[1247:1240] ,data[1255:1248] ,data[1263:1256] ,data[1271:1264] ,data[1279:1272] };
end
102 :begin
 dPIn = {data[359:352] ,data[367:360] ,data[375:368] ,data[383:376] ,data[391:384] ,data[583:576] ,data[591:584] ,data[599:592] ,data[607:600] ,data[615:608] ,data[807:800] ,data[815:808] ,data[823:816] ,data[831:824] ,data[839:832] ,data[1031:1024] ,data[1039:1032] ,data[1047:1040] ,data[1055:1048] ,data[1063:1056] ,data[1255:1248] ,data[1263:1256] ,data[1271:1264] ,data[1279:1272] ,data[1287:1280] };
end
103 :begin
 dPIn = {data[367:360] ,data[375:368] ,data[383:376] ,data[391:384] ,data[399:392] ,data[591:584] ,data[599:592] ,data[607:600] ,data[615:608] ,data[623:616] ,data[815:808] ,data[823:816] ,data[831:824] ,data[839:832] ,data[847:840] ,data[1039:1032] ,data[1047:1040] ,data[1055:1048] ,data[1063:1056] ,data[1071:1064] ,data[1263:1256] ,data[1271:1264] ,data[1279:1272] ,data[1287:1280] ,data[1295:1288] };
end
104 :begin
 dPIn = {data[375:368] ,data[383:376] ,data[391:384] ,data[399:392] ,data[407:400] ,data[599:592] ,data[607:600] ,data[615:608] ,data[623:616] ,data[631:624] ,data[823:816] ,data[831:824] ,data[839:832] ,data[847:840] ,data[855:848] ,data[1047:1040] ,data[1055:1048] ,data[1063:1056] ,data[1071:1064] ,data[1079:1072] ,data[1271:1264] ,data[1279:1272] ,data[1287:1280] ,data[1295:1288] ,data[1303:1296] };
end
105 :begin
 dPIn = {data[383:376] ,data[391:384] ,data[399:392] ,data[407:400] ,data[415:408] ,data[607:600] ,data[615:608] ,data[623:616] ,data[631:624] ,data[639:632] ,data[831:824] ,data[839:832] ,data[847:840] ,data[855:848] ,data[863:856] ,data[1055:1048] ,data[1063:1056] ,data[1071:1064] ,data[1079:1072] ,data[1087:1080] ,data[1279:1272] ,data[1287:1280] ,data[1295:1288] ,data[1303:1296] ,data[1311:1304] };
end
106 :begin
 dPIn = {data[391:384] ,data[399:392] ,data[407:400] ,data[415:408] ,data[423:416] ,data[615:608] ,data[623:616] ,data[631:624] ,data[639:632] ,data[647:640] ,data[839:832] ,data[847:840] ,data[855:848] ,data[863:856] ,data[871:864] ,data[1063:1056] ,data[1071:1064] ,data[1079:1072] ,data[1087:1080] ,data[1095:1088] ,data[1287:1280] ,data[1295:1288] ,data[1303:1296] ,data[1311:1304] ,data[1319:1312] };
end
107 :begin
 dPIn = {data[399:392] ,data[407:400] ,data[415:408] ,data[423:416] ,data[431:424] ,data[623:616] ,data[631:624] ,data[639:632] ,data[647:640] ,data[655:648] ,data[847:840] ,data[855:848] ,data[863:856] ,data[871:864] ,data[879:872] ,data[1071:1064] ,data[1079:1072] ,data[1087:1080] ,data[1095:1088] ,data[1103:1096] ,data[1295:1288] ,data[1303:1296] ,data[1311:1304] ,data[1319:1312] ,data[1327:1320] };
end
108 :begin
 dPIn = {data[407:400] ,data[415:408] ,data[423:416] ,data[431:424] ,data[439:432] ,data[631:624] ,data[639:632] ,data[647:640] ,data[655:648] ,data[663:656] ,data[855:848] ,data[863:856] ,data[871:864] ,data[879:872] ,data[887:880] ,data[1079:1072] ,data[1087:1080] ,data[1095:1088] ,data[1103:1096] ,data[1111:1104] ,data[1303:1296] ,data[1311:1304] ,data[1319:1312] ,data[1327:1320] ,data[1335:1328] };
end
109 :begin
 dPIn = {data[415:408] ,data[423:416] ,data[431:424] ,data[439:432] ,data[447:440] ,data[639:632] ,data[647:640] ,data[655:648] ,data[663:656] ,data[671:664] ,data[863:856] ,data[871:864] ,data[879:872] ,data[887:880] ,data[895:888] ,data[1087:1080] ,data[1095:1088] ,data[1103:1096] ,data[1111:1104] ,data[1119:1112] ,data[1311:1304] ,data[1319:1312] ,data[1327:1320] ,data[1335:1328] ,data[1343:1336] };
end
110 :begin
 dPIn = {data[423:416] ,data[431:424] ,data[439:432] ,data[447:440] ,0 ,data[647:640] ,data[655:648] ,data[663:656] ,data[671:664] ,0 ,data[871:864] ,data[879:872] ,data[887:880] ,data[895:888] ,0 ,data[1095:1088] ,data[1103:1096] ,data[1111:1104] ,data[1119:1112] ,0 ,data[1319:1312] ,data[1327:1320] ,data[1335:1328] ,data[1343:1336] ,0 };
end
111 :begin
 dPIn = {data[431:424] ,data[439:432] ,data[447:440] ,0 ,0 ,data[655:648] ,data[663:656] ,data[671:664] ,0 ,0 ,data[879:872] ,data[887:880] ,data[895:888] ,0 ,0 ,data[1103:1096] ,data[1111:1104] ,data[1119:1112] ,0 ,0 ,data[1327:1320] ,data[1335:1328] ,data[1343:1336] ,0 ,0 };
end
112 :begin
 dPIn = {0 ,0 ,data[455:448] ,data[463:456] ,data[471:464] ,0 ,0 ,data[679:672] ,data[687:680] ,data[695:688] ,0 ,0 ,data[903:896] ,data[911:904] ,data[919:912] ,0 ,0 ,data[1127:1120] ,data[1135:1128] ,data[1143:1136] ,0 ,0 ,data[1351:1344] ,data[1359:1352] ,data[1367:1360] };
end
113 :begin
 dPIn = {0 ,data[455:448] ,data[463:456] ,data[471:464] ,data[479:472] ,0 ,data[679:672] ,data[687:680] ,data[695:688] ,data[703:696] ,0 ,data[903:896] ,data[911:904] ,data[919:912] ,data[927:920] ,0 ,data[1127:1120] ,data[1135:1128] ,data[1143:1136] ,data[1151:1144] ,0 ,data[1351:1344] ,data[1359:1352] ,data[1367:1360] ,data[1375:1368] };
end
114 :begin
 dPIn = {data[455:448] ,data[463:456] ,data[471:464] ,data[479:472] ,data[487:480] ,data[679:672] ,data[687:680] ,data[695:688] ,data[703:696] ,data[711:704] ,data[903:896] ,data[911:904] ,data[919:912] ,data[927:920] ,data[935:928] ,data[1127:1120] ,data[1135:1128] ,data[1143:1136] ,data[1151:1144] ,data[1159:1152] ,data[1351:1344] ,data[1359:1352] ,data[1367:1360] ,data[1375:1368] ,data[1383:1376] };
end
115 :begin
 dPIn = {data[463:456] ,data[471:464] ,data[479:472] ,data[487:480] ,data[495:488] ,data[687:680] ,data[695:688] ,data[703:696] ,data[711:704] ,data[719:712] ,data[911:904] ,data[919:912] ,data[927:920] ,data[935:928] ,data[943:936] ,data[1135:1128] ,data[1143:1136] ,data[1151:1144] ,data[1159:1152] ,data[1167:1160] ,data[1359:1352] ,data[1367:1360] ,data[1375:1368] ,data[1383:1376] ,data[1391:1384] };
end
116 :begin
 dPIn = {data[471:464] ,data[479:472] ,data[487:480] ,data[495:488] ,data[503:496] ,data[695:688] ,data[703:696] ,data[711:704] ,data[719:712] ,data[727:720] ,data[919:912] ,data[927:920] ,data[935:928] ,data[943:936] ,data[951:944] ,data[1143:1136] ,data[1151:1144] ,data[1159:1152] ,data[1167:1160] ,data[1175:1168] ,data[1367:1360] ,data[1375:1368] ,data[1383:1376] ,data[1391:1384] ,data[1399:1392] };
end
117 :begin
 dPIn = {data[479:472] ,data[487:480] ,data[495:488] ,data[503:496] ,data[511:504] ,data[703:696] ,data[711:704] ,data[719:712] ,data[727:720] ,data[735:728] ,data[927:920] ,data[935:928] ,data[943:936] ,data[951:944] ,data[959:952] ,data[1151:1144] ,data[1159:1152] ,data[1167:1160] ,data[1175:1168] ,data[1183:1176] ,data[1375:1368] ,data[1383:1376] ,data[1391:1384] ,data[1399:1392] ,data[1407:1400] };
end
118 :begin
 dPIn = {data[487:480] ,data[495:488] ,data[503:496] ,data[511:504] ,data[519:512] ,data[711:704] ,data[719:712] ,data[727:720] ,data[735:728] ,data[743:736] ,data[935:928] ,data[943:936] ,data[951:944] ,data[959:952] ,data[967:960] ,data[1159:1152] ,data[1167:1160] ,data[1175:1168] ,data[1183:1176] ,data[1191:1184] ,data[1383:1376] ,data[1391:1384] ,data[1399:1392] ,data[1407:1400] ,data[1415:1408] };
end
119 :begin
 dPIn = {data[495:488] ,data[503:496] ,data[511:504] ,data[519:512] ,data[527:520] ,data[719:712] ,data[727:720] ,data[735:728] ,data[743:736] ,data[751:744] ,data[943:936] ,data[951:944] ,data[959:952] ,data[967:960] ,data[975:968] ,data[1167:1160] ,data[1175:1168] ,data[1183:1176] ,data[1191:1184] ,data[1199:1192] ,data[1391:1384] ,data[1399:1392] ,data[1407:1400] ,data[1415:1408] ,data[1423:1416] };
end
120 :begin
 dPIn = {data[503:496] ,data[511:504] ,data[519:512] ,data[527:520] ,data[535:528] ,data[727:720] ,data[735:728] ,data[743:736] ,data[751:744] ,data[759:752] ,data[951:944] ,data[959:952] ,data[967:960] ,data[975:968] ,data[983:976] ,data[1175:1168] ,data[1183:1176] ,data[1191:1184] ,data[1199:1192] ,data[1207:1200] ,data[1399:1392] ,data[1407:1400] ,data[1415:1408] ,data[1423:1416] ,data[1431:1424] };
end
121 :begin
 dPIn = {data[511:504] ,data[519:512] ,data[527:520] ,data[535:528] ,data[543:536] ,data[735:728] ,data[743:736] ,data[751:744] ,data[759:752] ,data[767:760] ,data[959:952] ,data[967:960] ,data[975:968] ,data[983:976] ,data[991:984] ,data[1183:1176] ,data[1191:1184] ,data[1199:1192] ,data[1207:1200] ,data[1215:1208] ,data[1407:1400] ,data[1415:1408] ,data[1423:1416] ,data[1431:1424] ,data[1439:1432] };
end
122 :begin
 dPIn = {data[519:512] ,data[527:520] ,data[535:528] ,data[543:536] ,data[551:544] ,data[743:736] ,data[751:744] ,data[759:752] ,data[767:760] ,data[775:768] ,data[967:960] ,data[975:968] ,data[983:976] ,data[991:984] ,data[999:992] ,data[1191:1184] ,data[1199:1192] ,data[1207:1200] ,data[1215:1208] ,data[1223:1216] ,data[1415:1408] ,data[1423:1416] ,data[1431:1424] ,data[1439:1432] ,data[1447:1440] };
end
123 :begin
 dPIn = {data[527:520] ,data[535:528] ,data[543:536] ,data[551:544] ,data[559:552] ,data[751:744] ,data[759:752] ,data[767:760] ,data[775:768] ,data[783:776] ,data[975:968] ,data[983:976] ,data[991:984] ,data[999:992] ,data[1007:1000] ,data[1199:1192] ,data[1207:1200] ,data[1215:1208] ,data[1223:1216] ,data[1231:1224] ,data[1423:1416] ,data[1431:1424] ,data[1439:1432] ,data[1447:1440] ,data[1455:1448] };
end
124 :begin
 dPIn = {data[535:528] ,data[543:536] ,data[551:544] ,data[559:552] ,data[567:560] ,data[759:752] ,data[767:760] ,data[775:768] ,data[783:776] ,data[791:784] ,data[983:976] ,data[991:984] ,data[999:992] ,data[1007:1000] ,data[1015:1008] ,data[1207:1200] ,data[1215:1208] ,data[1223:1216] ,data[1231:1224] ,data[1239:1232] ,data[1431:1424] ,data[1439:1432] ,data[1447:1440] ,data[1455:1448] ,data[1463:1456] };
end
125 :begin
 dPIn = {data[543:536] ,data[551:544] ,data[559:552] ,data[567:560] ,data[575:568] ,data[767:760] ,data[775:768] ,data[783:776] ,data[791:784] ,data[799:792] ,data[991:984] ,data[999:992] ,data[1007:1000] ,data[1015:1008] ,data[1023:1016] ,data[1215:1208] ,data[1223:1216] ,data[1231:1224] ,data[1239:1232] ,data[1247:1240] ,data[1439:1432] ,data[1447:1440] ,data[1455:1448] ,data[1463:1456] ,data[1471:1464] };
end
126 :begin
 dPIn = {data[551:544] ,data[559:552] ,data[567:560] ,data[575:568] ,data[583:576] ,data[775:768] ,data[783:776] ,data[791:784] ,data[799:792] ,data[807:800] ,data[999:992] ,data[1007:1000] ,data[1015:1008] ,data[1023:1016] ,data[1031:1024] ,data[1223:1216] ,data[1231:1224] ,data[1239:1232] ,data[1247:1240] ,data[1255:1248] ,data[1447:1440] ,data[1455:1448] ,data[1463:1456] ,data[1471:1464] ,data[1479:1472] };
end
127 :begin
 dPIn = {data[559:552] ,data[567:560] ,data[575:568] ,data[583:576] ,data[591:584] ,data[783:776] ,data[791:784] ,data[799:792] ,data[807:800] ,data[815:808] ,data[1007:1000] ,data[1015:1008] ,data[1023:1016] ,data[1031:1024] ,data[1039:1032] ,data[1231:1224] ,data[1239:1232] ,data[1247:1240] ,data[1255:1248] ,data[1263:1256] ,data[1455:1448] ,data[1463:1456] ,data[1471:1464] ,data[1479:1472] ,data[1487:1480] };
end
128 :begin
 dPIn = {data[567:560] ,data[575:568] ,data[583:576] ,data[591:584] ,data[599:592] ,data[791:784] ,data[799:792] ,data[807:800] ,data[815:808] ,data[823:816] ,data[1015:1008] ,data[1023:1016] ,data[1031:1024] ,data[1039:1032] ,data[1047:1040] ,data[1239:1232] ,data[1247:1240] ,data[1255:1248] ,data[1263:1256] ,data[1271:1264] ,data[1463:1456] ,data[1471:1464] ,data[1479:1472] ,data[1487:1480] ,data[1495:1488] };
end
129 :begin
 dPIn = {data[575:568] ,data[583:576] ,data[591:584] ,data[599:592] ,data[607:600] ,data[799:792] ,data[807:800] ,data[815:808] ,data[823:816] ,data[831:824] ,data[1023:1016] ,data[1031:1024] ,data[1039:1032] ,data[1047:1040] ,data[1055:1048] ,data[1247:1240] ,data[1255:1248] ,data[1263:1256] ,data[1271:1264] ,data[1279:1272] ,data[1471:1464] ,data[1479:1472] ,data[1487:1480] ,data[1495:1488] ,data[1503:1496] };
end
130 :begin
 dPIn = {data[583:576] ,data[591:584] ,data[599:592] ,data[607:600] ,data[615:608] ,data[807:800] ,data[815:808] ,data[823:816] ,data[831:824] ,data[839:832] ,data[1031:1024] ,data[1039:1032] ,data[1047:1040] ,data[1055:1048] ,data[1063:1056] ,data[1255:1248] ,data[1263:1256] ,data[1271:1264] ,data[1279:1272] ,data[1287:1280] ,data[1479:1472] ,data[1487:1480] ,data[1495:1488] ,data[1503:1496] ,data[1511:1504] };
end
131 :begin
 dPIn = {data[591:584] ,data[599:592] ,data[607:600] ,data[615:608] ,data[623:616] ,data[815:808] ,data[823:816] ,data[831:824] ,data[839:832] ,data[847:840] ,data[1039:1032] ,data[1047:1040] ,data[1055:1048] ,data[1063:1056] ,data[1071:1064] ,data[1263:1256] ,data[1271:1264] ,data[1279:1272] ,data[1287:1280] ,data[1295:1288] ,data[1487:1480] ,data[1495:1488] ,data[1503:1496] ,data[1511:1504] ,data[1519:1512] };
end
132 :begin
 dPIn = {data[599:592] ,data[607:600] ,data[615:608] ,data[623:616] ,data[631:624] ,data[823:816] ,data[831:824] ,data[839:832] ,data[847:840] ,data[855:848] ,data[1047:1040] ,data[1055:1048] ,data[1063:1056] ,data[1071:1064] ,data[1079:1072] ,data[1271:1264] ,data[1279:1272] ,data[1287:1280] ,data[1295:1288] ,data[1303:1296] ,data[1495:1488] ,data[1503:1496] ,data[1511:1504] ,data[1519:1512] ,data[1527:1520] };
end
133 :begin
 dPIn = {data[607:600] ,data[615:608] ,data[623:616] ,data[631:624] ,data[639:632] ,data[831:824] ,data[839:832] ,data[847:840] ,data[855:848] ,data[863:856] ,data[1055:1048] ,data[1063:1056] ,data[1071:1064] ,data[1079:1072] ,data[1087:1080] ,data[1279:1272] ,data[1287:1280] ,data[1295:1288] ,data[1303:1296] ,data[1311:1304] ,data[1503:1496] ,data[1511:1504] ,data[1519:1512] ,data[1527:1520] ,data[1535:1528] };
end
134 :begin
 dPIn = {data[615:608] ,data[623:616] ,data[631:624] ,data[639:632] ,data[647:640] ,data[839:832] ,data[847:840] ,data[855:848] ,data[863:856] ,data[871:864] ,data[1063:1056] ,data[1071:1064] ,data[1079:1072] ,data[1087:1080] ,data[1095:1088] ,data[1287:1280] ,data[1295:1288] ,data[1303:1296] ,data[1311:1304] ,data[1319:1312] ,data[1511:1504] ,data[1519:1512] ,data[1527:1520] ,data[1535:1528] ,data[1543:1536] };
end
135 :begin
 dPIn = {data[623:616] ,data[631:624] ,data[639:632] ,data[647:640] ,data[655:648] ,data[847:840] ,data[855:848] ,data[863:856] ,data[871:864] ,data[879:872] ,data[1071:1064] ,data[1079:1072] ,data[1087:1080] ,data[1095:1088] ,data[1103:1096] ,data[1295:1288] ,data[1303:1296] ,data[1311:1304] ,data[1319:1312] ,data[1327:1320] ,data[1519:1512] ,data[1527:1520] ,data[1535:1528] ,data[1543:1536] ,data[1551:1544] };
end
136 :begin
 dPIn = {data[631:624] ,data[639:632] ,data[647:640] ,data[655:648] ,data[663:656] ,data[855:848] ,data[863:856] ,data[871:864] ,data[879:872] ,data[887:880] ,data[1079:1072] ,data[1087:1080] ,data[1095:1088] ,data[1103:1096] ,data[1111:1104] ,data[1303:1296] ,data[1311:1304] ,data[1319:1312] ,data[1327:1320] ,data[1335:1328] ,data[1527:1520] ,data[1535:1528] ,data[1543:1536] ,data[1551:1544] ,data[1559:1552] };
end
137 :begin
 dPIn = {data[639:632] ,data[647:640] ,data[655:648] ,data[663:656] ,data[671:664] ,data[863:856] ,data[871:864] ,data[879:872] ,data[887:880] ,data[895:888] ,data[1087:1080] ,data[1095:1088] ,data[1103:1096] ,data[1111:1104] ,data[1119:1112] ,data[1311:1304] ,data[1319:1312] ,data[1327:1320] ,data[1335:1328] ,data[1343:1336] ,data[1535:1528] ,data[1543:1536] ,data[1551:1544] ,data[1559:1552] ,data[1567:1560] };
end
138 :begin
 dPIn = {data[647:640] ,data[655:648] ,data[663:656] ,data[671:664] ,0 ,data[871:864] ,data[879:872] ,data[887:880] ,data[895:888] ,0 ,data[1095:1088] ,data[1103:1096] ,data[1111:1104] ,data[1119:1112] ,0 ,data[1319:1312] ,data[1327:1320] ,data[1335:1328] ,data[1343:1336] ,0 ,data[1543:1536] ,data[1551:1544] ,data[1559:1552] ,data[1567:1560] ,0 };
end
139 :begin
 dPIn = {data[655:648] ,data[663:656] ,data[671:664] ,0 ,0 ,data[879:872] ,data[887:880] ,data[895:888] ,0 ,0 ,data[1103:1096] ,data[1111:1104] ,data[1119:1112] ,0 ,0 ,data[1327:1320] ,data[1335:1328] ,data[1343:1336] ,0 ,0 ,data[1551:1544] ,data[1559:1552] ,data[1567:1560] ,0 ,0 };
end
140 :begin
 dPIn = {0 ,0 ,data[679:672] ,data[687:680] ,data[695:688] ,0 ,0 ,data[903:896] ,data[911:904] ,data[919:912] ,0 ,0 ,data[1127:1120] ,data[1135:1128] ,data[1143:1136] ,0 ,0 ,data[1351:1344] ,data[1359:1352] ,data[1367:1360] ,0 ,0 ,data[1575:1568] ,data[1583:1576] ,data[1591:1584] };
end
141 :begin
 dPIn = {0 ,data[679:672] ,data[687:680] ,data[695:688] ,data[703:696] ,0 ,data[903:896] ,data[911:904] ,data[919:912] ,data[927:920] ,0 ,data[1127:1120] ,data[1135:1128] ,data[1143:1136] ,data[1151:1144] ,0 ,data[1351:1344] ,data[1359:1352] ,data[1367:1360] ,data[1375:1368] ,0 ,data[1575:1568] ,data[1583:1576] ,data[1591:1584] ,data[1599:1592] };
end
142 :begin
 dPIn = {data[679:672] ,data[687:680] ,data[695:688] ,data[703:696] ,data[711:704] ,data[903:896] ,data[911:904] ,data[919:912] ,data[927:920] ,data[935:928] ,data[1127:1120] ,data[1135:1128] ,data[1143:1136] ,data[1151:1144] ,data[1159:1152] ,data[1351:1344] ,data[1359:1352] ,data[1367:1360] ,data[1375:1368] ,data[1383:1376] ,data[1575:1568] ,data[1583:1576] ,data[1591:1584] ,data[1599:1592] ,data[1607:1600] };
end
143 :begin
 dPIn = {data[687:680] ,data[695:688] ,data[703:696] ,data[711:704] ,data[719:712] ,data[911:904] ,data[919:912] ,data[927:920] ,data[935:928] ,data[943:936] ,data[1135:1128] ,data[1143:1136] ,data[1151:1144] ,data[1159:1152] ,data[1167:1160] ,data[1359:1352] ,data[1367:1360] ,data[1375:1368] ,data[1383:1376] ,data[1391:1384] ,data[1583:1576] ,data[1591:1584] ,data[1599:1592] ,data[1607:1600] ,data[1615:1608] };
end
144 :begin
 dPIn = {data[695:688] ,data[703:696] ,data[711:704] ,data[719:712] ,data[727:720] ,data[919:912] ,data[927:920] ,data[935:928] ,data[943:936] ,data[951:944] ,data[1143:1136] ,data[1151:1144] ,data[1159:1152] ,data[1167:1160] ,data[1175:1168] ,data[1367:1360] ,data[1375:1368] ,data[1383:1376] ,data[1391:1384] ,data[1399:1392] ,data[1591:1584] ,data[1599:1592] ,data[1607:1600] ,data[1615:1608] ,data[1623:1616] };
end
145 :begin
 dPIn = {data[703:696] ,data[711:704] ,data[719:712] ,data[727:720] ,data[735:728] ,data[927:920] ,data[935:928] ,data[943:936] ,data[951:944] ,data[959:952] ,data[1151:1144] ,data[1159:1152] ,data[1167:1160] ,data[1175:1168] ,data[1183:1176] ,data[1375:1368] ,data[1383:1376] ,data[1391:1384] ,data[1399:1392] ,data[1407:1400] ,data[1599:1592] ,data[1607:1600] ,data[1615:1608] ,data[1623:1616] ,data[1631:1624] };
end
146 :begin
 dPIn = {data[711:704] ,data[719:712] ,data[727:720] ,data[735:728] ,data[743:736] ,data[935:928] ,data[943:936] ,data[951:944] ,data[959:952] ,data[967:960] ,data[1159:1152] ,data[1167:1160] ,data[1175:1168] ,data[1183:1176] ,data[1191:1184] ,data[1383:1376] ,data[1391:1384] ,data[1399:1392] ,data[1407:1400] ,data[1415:1408] ,data[1607:1600] ,data[1615:1608] ,data[1623:1616] ,data[1631:1624] ,data[1639:1632] };
end
147 :begin
 dPIn = {data[719:712] ,data[727:720] ,data[735:728] ,data[743:736] ,data[751:744] ,data[943:936] ,data[951:944] ,data[959:952] ,data[967:960] ,data[975:968] ,data[1167:1160] ,data[1175:1168] ,data[1183:1176] ,data[1191:1184] ,data[1199:1192] ,data[1391:1384] ,data[1399:1392] ,data[1407:1400] ,data[1415:1408] ,data[1423:1416] ,data[1615:1608] ,data[1623:1616] ,data[1631:1624] ,data[1639:1632] ,data[1647:1640] };
end
148 :begin
 dPIn = {data[727:720] ,data[735:728] ,data[743:736] ,data[751:744] ,data[759:752] ,data[951:944] ,data[959:952] ,data[967:960] ,data[975:968] ,data[983:976] ,data[1175:1168] ,data[1183:1176] ,data[1191:1184] ,data[1199:1192] ,data[1207:1200] ,data[1399:1392] ,data[1407:1400] ,data[1415:1408] ,data[1423:1416] ,data[1431:1424] ,data[1623:1616] ,data[1631:1624] ,data[1639:1632] ,data[1647:1640] ,data[1655:1648] };
end
149 :begin
 dPIn = {data[735:728] ,data[743:736] ,data[751:744] ,data[759:752] ,data[767:760] ,data[959:952] ,data[967:960] ,data[975:968] ,data[983:976] ,data[991:984] ,data[1183:1176] ,data[1191:1184] ,data[1199:1192] ,data[1207:1200] ,data[1215:1208] ,data[1407:1400] ,data[1415:1408] ,data[1423:1416] ,data[1431:1424] ,data[1439:1432] ,data[1631:1624] ,data[1639:1632] ,data[1647:1640] ,data[1655:1648] ,data[1663:1656] };
end
150 :begin
 dPIn = {data[743:736] ,data[751:744] ,data[759:752] ,data[767:760] ,data[775:768] ,data[967:960] ,data[975:968] ,data[983:976] ,data[991:984] ,data[999:992] ,data[1191:1184] ,data[1199:1192] ,data[1207:1200] ,data[1215:1208] ,data[1223:1216] ,data[1415:1408] ,data[1423:1416] ,data[1431:1424] ,data[1439:1432] ,data[1447:1440] ,data[1639:1632] ,data[1647:1640] ,data[1655:1648] ,data[1663:1656] ,data[1671:1664] };
end
151 :begin
 dPIn = {data[751:744] ,data[759:752] ,data[767:760] ,data[775:768] ,data[783:776] ,data[975:968] ,data[983:976] ,data[991:984] ,data[999:992] ,data[1007:1000] ,data[1199:1192] ,data[1207:1200] ,data[1215:1208] ,data[1223:1216] ,data[1231:1224] ,data[1423:1416] ,data[1431:1424] ,data[1439:1432] ,data[1447:1440] ,data[1455:1448] ,data[1647:1640] ,data[1655:1648] ,data[1663:1656] ,data[1671:1664] ,data[1679:1672] };
end
152 :begin
 dPIn = {data[759:752] ,data[767:760] ,data[775:768] ,data[783:776] ,data[791:784] ,data[983:976] ,data[991:984] ,data[999:992] ,data[1007:1000] ,data[1015:1008] ,data[1207:1200] ,data[1215:1208] ,data[1223:1216] ,data[1231:1224] ,data[1239:1232] ,data[1431:1424] ,data[1439:1432] ,data[1447:1440] ,data[1455:1448] ,data[1463:1456] ,data[1655:1648] ,data[1663:1656] ,data[1671:1664] ,data[1679:1672] ,data[1687:1680] };
end
153 :begin
 dPIn = {data[767:760] ,data[775:768] ,data[783:776] ,data[791:784] ,data[799:792] ,data[991:984] ,data[999:992] ,data[1007:1000] ,data[1015:1008] ,data[1023:1016] ,data[1215:1208] ,data[1223:1216] ,data[1231:1224] ,data[1239:1232] ,data[1247:1240] ,data[1439:1432] ,data[1447:1440] ,data[1455:1448] ,data[1463:1456] ,data[1471:1464] ,data[1663:1656] ,data[1671:1664] ,data[1679:1672] ,data[1687:1680] ,data[1695:1688] };
end
154 :begin
 dPIn = {data[775:768] ,data[783:776] ,data[791:784] ,data[799:792] ,data[807:800] ,data[999:992] ,data[1007:1000] ,data[1015:1008] ,data[1023:1016] ,data[1031:1024] ,data[1223:1216] ,data[1231:1224] ,data[1239:1232] ,data[1247:1240] ,data[1255:1248] ,data[1447:1440] ,data[1455:1448] ,data[1463:1456] ,data[1471:1464] ,data[1479:1472] ,data[1671:1664] ,data[1679:1672] ,data[1687:1680] ,data[1695:1688] ,data[1703:1696] };
end
155 :begin
 dPIn = {data[783:776] ,data[791:784] ,data[799:792] ,data[807:800] ,data[815:808] ,data[1007:1000] ,data[1015:1008] ,data[1023:1016] ,data[1031:1024] ,data[1039:1032] ,data[1231:1224] ,data[1239:1232] ,data[1247:1240] ,data[1255:1248] ,data[1263:1256] ,data[1455:1448] ,data[1463:1456] ,data[1471:1464] ,data[1479:1472] ,data[1487:1480] ,data[1679:1672] ,data[1687:1680] ,data[1695:1688] ,data[1703:1696] ,data[1711:1704] };
end
156 :begin
 dPIn = {data[791:784] ,data[799:792] ,data[807:800] ,data[815:808] ,data[823:816] ,data[1015:1008] ,data[1023:1016] ,data[1031:1024] ,data[1039:1032] ,data[1047:1040] ,data[1239:1232] ,data[1247:1240] ,data[1255:1248] ,data[1263:1256] ,data[1271:1264] ,data[1463:1456] ,data[1471:1464] ,data[1479:1472] ,data[1487:1480] ,data[1495:1488] ,data[1687:1680] ,data[1695:1688] ,data[1703:1696] ,data[1711:1704] ,data[1719:1712] };
end
157 :begin
 dPIn = {data[799:792] ,data[807:800] ,data[815:808] ,data[823:816] ,data[831:824] ,data[1023:1016] ,data[1031:1024] ,data[1039:1032] ,data[1047:1040] ,data[1055:1048] ,data[1247:1240] ,data[1255:1248] ,data[1263:1256] ,data[1271:1264] ,data[1279:1272] ,data[1471:1464] ,data[1479:1472] ,data[1487:1480] ,data[1495:1488] ,data[1503:1496] ,data[1695:1688] ,data[1703:1696] ,data[1711:1704] ,data[1719:1712] ,data[1727:1720] };
end
158 :begin
 dPIn = {data[807:800] ,data[815:808] ,data[823:816] ,data[831:824] ,data[839:832] ,data[1031:1024] ,data[1039:1032] ,data[1047:1040] ,data[1055:1048] ,data[1063:1056] ,data[1255:1248] ,data[1263:1256] ,data[1271:1264] ,data[1279:1272] ,data[1287:1280] ,data[1479:1472] ,data[1487:1480] ,data[1495:1488] ,data[1503:1496] ,data[1511:1504] ,data[1703:1696] ,data[1711:1704] ,data[1719:1712] ,data[1727:1720] ,data[1735:1728] };
end
159 :begin
 dPIn = {data[815:808] ,data[823:816] ,data[831:824] ,data[839:832] ,data[847:840] ,data[1039:1032] ,data[1047:1040] ,data[1055:1048] ,data[1063:1056] ,data[1071:1064] ,data[1263:1256] ,data[1271:1264] ,data[1279:1272] ,data[1287:1280] ,data[1295:1288] ,data[1487:1480] ,data[1495:1488] ,data[1503:1496] ,data[1511:1504] ,data[1519:1512] ,data[1711:1704] ,data[1719:1712] ,data[1727:1720] ,data[1735:1728] ,data[1743:1736] };
end
160 :begin
 dPIn = {data[823:816] ,data[831:824] ,data[839:832] ,data[847:840] ,data[855:848] ,data[1047:1040] ,data[1055:1048] ,data[1063:1056] ,data[1071:1064] ,data[1079:1072] ,data[1271:1264] ,data[1279:1272] ,data[1287:1280] ,data[1295:1288] ,data[1303:1296] ,data[1495:1488] ,data[1503:1496] ,data[1511:1504] ,data[1519:1512] ,data[1527:1520] ,data[1719:1712] ,data[1727:1720] ,data[1735:1728] ,data[1743:1736] ,data[1751:1744] };
end
161 :begin
 dPIn = {data[831:824] ,data[839:832] ,data[847:840] ,data[855:848] ,data[863:856] ,data[1055:1048] ,data[1063:1056] ,data[1071:1064] ,data[1079:1072] ,data[1087:1080] ,data[1279:1272] ,data[1287:1280] ,data[1295:1288] ,data[1303:1296] ,data[1311:1304] ,data[1503:1496] ,data[1511:1504] ,data[1519:1512] ,data[1527:1520] ,data[1535:1528] ,data[1727:1720] ,data[1735:1728] ,data[1743:1736] ,data[1751:1744] ,data[1759:1752] };
end
162 :begin
 dPIn = {data[839:832] ,data[847:840] ,data[855:848] ,data[863:856] ,data[871:864] ,data[1063:1056] ,data[1071:1064] ,data[1079:1072] ,data[1087:1080] ,data[1095:1088] ,data[1287:1280] ,data[1295:1288] ,data[1303:1296] ,data[1311:1304] ,data[1319:1312] ,data[1511:1504] ,data[1519:1512] ,data[1527:1520] ,data[1535:1528] ,data[1543:1536] ,data[1735:1728] ,data[1743:1736] ,data[1751:1744] ,data[1759:1752] ,data[1767:1760] };
end
163 :begin
 dPIn = {data[847:840] ,data[855:848] ,data[863:856] ,data[871:864] ,data[879:872] ,data[1071:1064] ,data[1079:1072] ,data[1087:1080] ,data[1095:1088] ,data[1103:1096] ,data[1295:1288] ,data[1303:1296] ,data[1311:1304] ,data[1319:1312] ,data[1327:1320] ,data[1519:1512] ,data[1527:1520] ,data[1535:1528] ,data[1543:1536] ,data[1551:1544] ,data[1743:1736] ,data[1751:1744] ,data[1759:1752] ,data[1767:1760] ,data[1775:1768] };
end
164 :begin
 dPIn = {data[855:848] ,data[863:856] ,data[871:864] ,data[879:872] ,data[887:880] ,data[1079:1072] ,data[1087:1080] ,data[1095:1088] ,data[1103:1096] ,data[1111:1104] ,data[1303:1296] ,data[1311:1304] ,data[1319:1312] ,data[1327:1320] ,data[1335:1328] ,data[1527:1520] ,data[1535:1528] ,data[1543:1536] ,data[1551:1544] ,data[1559:1552] ,data[1751:1744] ,data[1759:1752] ,data[1767:1760] ,data[1775:1768] ,data[1783:1776] };
end
165 :begin
 dPIn = {data[863:856] ,data[871:864] ,data[879:872] ,data[887:880] ,data[895:888] ,data[1087:1080] ,data[1095:1088] ,data[1103:1096] ,data[1111:1104] ,data[1119:1112] ,data[1311:1304] ,data[1319:1312] ,data[1327:1320] ,data[1335:1328] ,data[1343:1336] ,data[1535:1528] ,data[1543:1536] ,data[1551:1544] ,data[1559:1552] ,data[1567:1560] ,data[1759:1752] ,data[1767:1760] ,data[1775:1768] ,data[1783:1776] ,data[1791:1784] };
end
166 :begin
 dPIn = {data[871:864] ,data[879:872] ,data[887:880] ,data[895:888] ,0 ,data[1095:1088] ,data[1103:1096] ,data[1111:1104] ,data[1119:1112] ,0 ,data[1319:1312] ,data[1327:1320] ,data[1335:1328] ,data[1343:1336] ,0 ,data[1543:1536] ,data[1551:1544] ,data[1559:1552] ,data[1567:1560] ,0 ,data[1767:1760] ,data[1775:1768] ,data[1783:1776] ,data[1791:1784] ,0 };
end
167 :begin
 dPIn = {data[879:872] ,data[887:880] ,data[895:888] ,0 ,0 ,data[1103:1096] ,data[1111:1104] ,data[1119:1112] ,0 ,0 ,data[1327:1320] ,data[1335:1328] ,data[1343:1336] ,0 ,0 ,data[1551:1544] ,data[1559:1552] ,data[1567:1560] ,0 ,0 ,data[1775:1768] ,data[1783:1776] ,data[1791:1784] ,0 ,0 };
end
168 :begin
 dPIn = {0 ,0 ,data[903:896] ,data[911:904] ,data[919:912] ,0 ,0 ,data[1127:1120] ,data[1135:1128] ,data[1143:1136] ,0 ,0 ,data[1351:1344] ,data[1359:1352] ,data[1367:1360] ,0 ,0 ,data[1575:1568] ,data[1583:1576] ,data[1591:1584] ,0 ,0 ,data[1799:1792] ,data[1807:1800] ,data[1815:1808] };
end
169 :begin
 dPIn = {0 ,data[903:896] ,data[911:904] ,data[919:912] ,data[927:920] ,0 ,data[1127:1120] ,data[1135:1128] ,data[1143:1136] ,data[1151:1144] ,0 ,data[1351:1344] ,data[1359:1352] ,data[1367:1360] ,data[1375:1368] ,0 ,data[1575:1568] ,data[1583:1576] ,data[1591:1584] ,data[1599:1592] ,0 ,data[1799:1792] ,data[1807:1800] ,data[1815:1808] ,data[1823:1816] };
end
170 :begin
 dPIn = {data[903:896] ,data[911:904] ,data[919:912] ,data[927:920] ,data[935:928] ,data[1127:1120] ,data[1135:1128] ,data[1143:1136] ,data[1151:1144] ,data[1159:1152] ,data[1351:1344] ,data[1359:1352] ,data[1367:1360] ,data[1375:1368] ,data[1383:1376] ,data[1575:1568] ,data[1583:1576] ,data[1591:1584] ,data[1599:1592] ,data[1607:1600] ,data[1799:1792] ,data[1807:1800] ,data[1815:1808] ,data[1823:1816] ,data[1831:1824] };
end
171 :begin
 dPIn = {data[911:904] ,data[919:912] ,data[927:920] ,data[935:928] ,data[943:936] ,data[1135:1128] ,data[1143:1136] ,data[1151:1144] ,data[1159:1152] ,data[1167:1160] ,data[1359:1352] ,data[1367:1360] ,data[1375:1368] ,data[1383:1376] ,data[1391:1384] ,data[1583:1576] ,data[1591:1584] ,data[1599:1592] ,data[1607:1600] ,data[1615:1608] ,data[1807:1800] ,data[1815:1808] ,data[1823:1816] ,data[1831:1824] ,data[1839:1832] };
end
172 :begin
 dPIn = {data[919:912] ,data[927:920] ,data[935:928] ,data[943:936] ,data[951:944] ,data[1143:1136] ,data[1151:1144] ,data[1159:1152] ,data[1167:1160] ,data[1175:1168] ,data[1367:1360] ,data[1375:1368] ,data[1383:1376] ,data[1391:1384] ,data[1399:1392] ,data[1591:1584] ,data[1599:1592] ,data[1607:1600] ,data[1615:1608] ,data[1623:1616] ,data[1815:1808] ,data[1823:1816] ,data[1831:1824] ,data[1839:1832] ,data[1847:1840] };
end
173 :begin
 dPIn = {data[927:920] ,data[935:928] ,data[943:936] ,data[951:944] ,data[959:952] ,data[1151:1144] ,data[1159:1152] ,data[1167:1160] ,data[1175:1168] ,data[1183:1176] ,data[1375:1368] ,data[1383:1376] ,data[1391:1384] ,data[1399:1392] ,data[1407:1400] ,data[1599:1592] ,data[1607:1600] ,data[1615:1608] ,data[1623:1616] ,data[1631:1624] ,data[1823:1816] ,data[1831:1824] ,data[1839:1832] ,data[1847:1840] ,data[1855:1848] };
end
174 :begin
 dPIn = {data[935:928] ,data[943:936] ,data[951:944] ,data[959:952] ,data[967:960] ,data[1159:1152] ,data[1167:1160] ,data[1175:1168] ,data[1183:1176] ,data[1191:1184] ,data[1383:1376] ,data[1391:1384] ,data[1399:1392] ,data[1407:1400] ,data[1415:1408] ,data[1607:1600] ,data[1615:1608] ,data[1623:1616] ,data[1631:1624] ,data[1639:1632] ,data[1831:1824] ,data[1839:1832] ,data[1847:1840] ,data[1855:1848] ,data[1863:1856] };
end
175 :begin
 dPIn = {data[943:936] ,data[951:944] ,data[959:952] ,data[967:960] ,data[975:968] ,data[1167:1160] ,data[1175:1168] ,data[1183:1176] ,data[1191:1184] ,data[1199:1192] ,data[1391:1384] ,data[1399:1392] ,data[1407:1400] ,data[1415:1408] ,data[1423:1416] ,data[1615:1608] ,data[1623:1616] ,data[1631:1624] ,data[1639:1632] ,data[1647:1640] ,data[1839:1832] ,data[1847:1840] ,data[1855:1848] ,data[1863:1856] ,data[1871:1864] };
end
176 :begin
 dPIn = {data[951:944] ,data[959:952] ,data[967:960] ,data[975:968] ,data[983:976] ,data[1175:1168] ,data[1183:1176] ,data[1191:1184] ,data[1199:1192] ,data[1207:1200] ,data[1399:1392] ,data[1407:1400] ,data[1415:1408] ,data[1423:1416] ,data[1431:1424] ,data[1623:1616] ,data[1631:1624] ,data[1639:1632] ,data[1647:1640] ,data[1655:1648] ,data[1847:1840] ,data[1855:1848] ,data[1863:1856] ,data[1871:1864] ,data[1879:1872] };
end
177 :begin
 dPIn = {data[959:952] ,data[967:960] ,data[975:968] ,data[983:976] ,data[991:984] ,data[1183:1176] ,data[1191:1184] ,data[1199:1192] ,data[1207:1200] ,data[1215:1208] ,data[1407:1400] ,data[1415:1408] ,data[1423:1416] ,data[1431:1424] ,data[1439:1432] ,data[1631:1624] ,data[1639:1632] ,data[1647:1640] ,data[1655:1648] ,data[1663:1656] ,data[1855:1848] ,data[1863:1856] ,data[1871:1864] ,data[1879:1872] ,data[1887:1880] };
end
178 :begin
 dPIn = {data[967:960] ,data[975:968] ,data[983:976] ,data[991:984] ,data[999:992] ,data[1191:1184] ,data[1199:1192] ,data[1207:1200] ,data[1215:1208] ,data[1223:1216] ,data[1415:1408] ,data[1423:1416] ,data[1431:1424] ,data[1439:1432] ,data[1447:1440] ,data[1639:1632] ,data[1647:1640] ,data[1655:1648] ,data[1663:1656] ,data[1671:1664] ,data[1863:1856] ,data[1871:1864] ,data[1879:1872] ,data[1887:1880] ,data[1895:1888] };
end
179 :begin
 dPIn = {data[975:968] ,data[983:976] ,data[991:984] ,data[999:992] ,data[1007:1000] ,data[1199:1192] ,data[1207:1200] ,data[1215:1208] ,data[1223:1216] ,data[1231:1224] ,data[1423:1416] ,data[1431:1424] ,data[1439:1432] ,data[1447:1440] ,data[1455:1448] ,data[1647:1640] ,data[1655:1648] ,data[1663:1656] ,data[1671:1664] ,data[1679:1672] ,data[1871:1864] ,data[1879:1872] ,data[1887:1880] ,data[1895:1888] ,data[1903:1896] };
end
180 :begin
 dPIn = {data[983:976] ,data[991:984] ,data[999:992] ,data[1007:1000] ,data[1015:1008] ,data[1207:1200] ,data[1215:1208] ,data[1223:1216] ,data[1231:1224] ,data[1239:1232] ,data[1431:1424] ,data[1439:1432] ,data[1447:1440] ,data[1455:1448] ,data[1463:1456] ,data[1655:1648] ,data[1663:1656] ,data[1671:1664] ,data[1679:1672] ,data[1687:1680] ,data[1879:1872] ,data[1887:1880] ,data[1895:1888] ,data[1903:1896] ,data[1911:1904] };
end
181 :begin
 dPIn = {data[991:984] ,data[999:992] ,data[1007:1000] ,data[1015:1008] ,data[1023:1016] ,data[1215:1208] ,data[1223:1216] ,data[1231:1224] ,data[1239:1232] ,data[1247:1240] ,data[1439:1432] ,data[1447:1440] ,data[1455:1448] ,data[1463:1456] ,data[1471:1464] ,data[1663:1656] ,data[1671:1664] ,data[1679:1672] ,data[1687:1680] ,data[1695:1688] ,data[1887:1880] ,data[1895:1888] ,data[1903:1896] ,data[1911:1904] ,data[1919:1912] };
end
182 :begin
 dPIn = {data[999:992] ,data[1007:1000] ,data[1015:1008] ,data[1023:1016] ,data[1031:1024] ,data[1223:1216] ,data[1231:1224] ,data[1239:1232] ,data[1247:1240] ,data[1255:1248] ,data[1447:1440] ,data[1455:1448] ,data[1463:1456] ,data[1471:1464] ,data[1479:1472] ,data[1671:1664] ,data[1679:1672] ,data[1687:1680] ,data[1695:1688] ,data[1703:1696] ,data[1895:1888] ,data[1903:1896] ,data[1911:1904] ,data[1919:1912] ,data[1927:1920] };
end
183 :begin
 dPIn = {data[1007:1000] ,data[1015:1008] ,data[1023:1016] ,data[1031:1024] ,data[1039:1032] ,data[1231:1224] ,data[1239:1232] ,data[1247:1240] ,data[1255:1248] ,data[1263:1256] ,data[1455:1448] ,data[1463:1456] ,data[1471:1464] ,data[1479:1472] ,data[1487:1480] ,data[1679:1672] ,data[1687:1680] ,data[1695:1688] ,data[1703:1696] ,data[1711:1704] ,data[1903:1896] ,data[1911:1904] ,data[1919:1912] ,data[1927:1920] ,data[1935:1928] };
end
184 :begin
 dPIn = {data[1015:1008] ,data[1023:1016] ,data[1031:1024] ,data[1039:1032] ,data[1047:1040] ,data[1239:1232] ,data[1247:1240] ,data[1255:1248] ,data[1263:1256] ,data[1271:1264] ,data[1463:1456] ,data[1471:1464] ,data[1479:1472] ,data[1487:1480] ,data[1495:1488] ,data[1687:1680] ,data[1695:1688] ,data[1703:1696] ,data[1711:1704] ,data[1719:1712] ,data[1911:1904] ,data[1919:1912] ,data[1927:1920] ,data[1935:1928] ,data[1943:1936] };
end
185 :begin
 dPIn = {data[1023:1016] ,data[1031:1024] ,data[1039:1032] ,data[1047:1040] ,data[1055:1048] ,data[1247:1240] ,data[1255:1248] ,data[1263:1256] ,data[1271:1264] ,data[1279:1272] ,data[1471:1464] ,data[1479:1472] ,data[1487:1480] ,data[1495:1488] ,data[1503:1496] ,data[1695:1688] ,data[1703:1696] ,data[1711:1704] ,data[1719:1712] ,data[1727:1720] ,data[1919:1912] ,data[1927:1920] ,data[1935:1928] ,data[1943:1936] ,data[1951:1944] };
end
186 :begin
 dPIn = {data[1031:1024] ,data[1039:1032] ,data[1047:1040] ,data[1055:1048] ,data[1063:1056] ,data[1255:1248] ,data[1263:1256] ,data[1271:1264] ,data[1279:1272] ,data[1287:1280] ,data[1479:1472] ,data[1487:1480] ,data[1495:1488] ,data[1503:1496] ,data[1511:1504] ,data[1703:1696] ,data[1711:1704] ,data[1719:1712] ,data[1727:1720] ,data[1735:1728] ,data[1927:1920] ,data[1935:1928] ,data[1943:1936] ,data[1951:1944] ,data[1959:1952] };
end
187 :begin
 dPIn = {data[1039:1032] ,data[1047:1040] ,data[1055:1048] ,data[1063:1056] ,data[1071:1064] ,data[1263:1256] ,data[1271:1264] ,data[1279:1272] ,data[1287:1280] ,data[1295:1288] ,data[1487:1480] ,data[1495:1488] ,data[1503:1496] ,data[1511:1504] ,data[1519:1512] ,data[1711:1704] ,data[1719:1712] ,data[1727:1720] ,data[1735:1728] ,data[1743:1736] ,data[1935:1928] ,data[1943:1936] ,data[1951:1944] ,data[1959:1952] ,data[1967:1960] };
end
188 :begin
 dPIn = {data[1047:1040] ,data[1055:1048] ,data[1063:1056] ,data[1071:1064] ,data[1079:1072] ,data[1271:1264] ,data[1279:1272] ,data[1287:1280] ,data[1295:1288] ,data[1303:1296] ,data[1495:1488] ,data[1503:1496] ,data[1511:1504] ,data[1519:1512] ,data[1527:1520] ,data[1719:1712] ,data[1727:1720] ,data[1735:1728] ,data[1743:1736] ,data[1751:1744] ,data[1943:1936] ,data[1951:1944] ,data[1959:1952] ,data[1967:1960] ,data[1975:1968] };
end
189 :begin
 dPIn = {data[1055:1048] ,data[1063:1056] ,data[1071:1064] ,data[1079:1072] ,data[1087:1080] ,data[1279:1272] ,data[1287:1280] ,data[1295:1288] ,data[1303:1296] ,data[1311:1304] ,data[1503:1496] ,data[1511:1504] ,data[1519:1512] ,data[1527:1520] ,data[1535:1528] ,data[1727:1720] ,data[1735:1728] ,data[1743:1736] ,data[1751:1744] ,data[1759:1752] ,data[1951:1944] ,data[1959:1952] ,data[1967:1960] ,data[1975:1968] ,data[1983:1976] };
end
190 :begin
 dPIn = {data[1063:1056] ,data[1071:1064] ,data[1079:1072] ,data[1087:1080] ,data[1095:1088] ,data[1287:1280] ,data[1295:1288] ,data[1303:1296] ,data[1311:1304] ,data[1319:1312] ,data[1511:1504] ,data[1519:1512] ,data[1527:1520] ,data[1535:1528] ,data[1543:1536] ,data[1735:1728] ,data[1743:1736] ,data[1751:1744] ,data[1759:1752] ,data[1767:1760] ,data[1959:1952] ,data[1967:1960] ,data[1975:1968] ,data[1983:1976] ,data[1991:1984] };
end
191 :begin
 dPIn = {data[1071:1064] ,data[1079:1072] ,data[1087:1080] ,data[1095:1088] ,data[1103:1096] ,data[1295:1288] ,data[1303:1296] ,data[1311:1304] ,data[1319:1312] ,data[1327:1320] ,data[1519:1512] ,data[1527:1520] ,data[1535:1528] ,data[1543:1536] ,data[1551:1544] ,data[1743:1736] ,data[1751:1744] ,data[1759:1752] ,data[1767:1760] ,data[1775:1768] ,data[1967:1960] ,data[1975:1968] ,data[1983:1976] ,data[1991:1984] ,data[1999:1992] };
end
192 :begin
 dPIn = {data[1079:1072] ,data[1087:1080] ,data[1095:1088] ,data[1103:1096] ,data[1111:1104] ,data[1303:1296] ,data[1311:1304] ,data[1319:1312] ,data[1327:1320] ,data[1335:1328] ,data[1527:1520] ,data[1535:1528] ,data[1543:1536] ,data[1551:1544] ,data[1559:1552] ,data[1751:1744] ,data[1759:1752] ,data[1767:1760] ,data[1775:1768] ,data[1783:1776] ,data[1975:1968] ,data[1983:1976] ,data[1991:1984] ,data[1999:1992] ,data[2007:2000] };
end
193 :begin
 dPIn = {data[1087:1080] ,data[1095:1088] ,data[1103:1096] ,data[1111:1104] ,data[1119:1112] ,data[1311:1304] ,data[1319:1312] ,data[1327:1320] ,data[1335:1328] ,data[1343:1336] ,data[1535:1528] ,data[1543:1536] ,data[1551:1544] ,data[1559:1552] ,data[1567:1560] ,data[1759:1752] ,data[1767:1760] ,data[1775:1768] ,data[1783:1776] ,data[1791:1784] ,data[1983:1976] ,data[1991:1984] ,data[1999:1992] ,data[2007:2000] ,data[2015:2008] };
end
194 :begin
 dPIn = {data[1095:1088] ,data[1103:1096] ,data[1111:1104] ,data[1119:1112] ,0 ,data[1319:1312] ,data[1327:1320] ,data[1335:1328] ,data[1343:1336] ,0 ,data[1543:1536] ,data[1551:1544] ,data[1559:1552] ,data[1567:1560] ,0 ,data[1767:1760] ,data[1775:1768] ,data[1783:1776] ,data[1791:1784] ,0 ,data[1991:1984] ,data[1999:1992] ,data[2007:2000] ,data[2015:2008] ,0 };
end
195 :begin
 dPIn = {data[1103:1096] ,data[1111:1104] ,data[1119:1112] ,0 ,0 ,data[1327:1320] ,data[1335:1328] ,data[1343:1336] ,0 ,0 ,data[1551:1544] ,data[1559:1552] ,data[1567:1560] ,0 ,0 ,data[1775:1768] ,data[1783:1776] ,data[1791:1784] ,0 ,0 ,data[1999:1992] ,data[2007:2000] ,data[2015:2008] ,0 ,0 };
end
196 :begin
 dPIn = {0 ,0 ,data[1127:1120] ,data[1135:1128] ,data[1143:1136] ,0 ,0 ,data[1351:1344] ,data[1359:1352] ,data[1367:1360] ,0 ,0 ,data[1575:1568] ,data[1583:1576] ,data[1591:1584] ,0 ,0 ,data[1799:1792] ,data[1807:1800] ,data[1815:1808] ,0 ,0 ,data[2023:2016] ,data[2031:2024] ,data[2039:2032] };
end
197 :begin
 dPIn = {0 ,data[1127:1120] ,data[1135:1128] ,data[1143:1136] ,data[1151:1144] ,0 ,data[1351:1344] ,data[1359:1352] ,data[1367:1360] ,data[1375:1368] ,0 ,data[1575:1568] ,data[1583:1576] ,data[1591:1584] ,data[1599:1592] ,0 ,data[1799:1792] ,data[1807:1800] ,data[1815:1808] ,data[1823:1816] ,0 ,data[2023:2016] ,data[2031:2024] ,data[2039:2032] ,data[2047:2040] };
end
198 :begin
 dPIn = {data[1127:1120] ,data[1135:1128] ,data[1143:1136] ,data[1151:1144] ,data[1159:1152] ,data[1351:1344] ,data[1359:1352] ,data[1367:1360] ,data[1375:1368] ,data[1383:1376] ,data[1575:1568] ,data[1583:1576] ,data[1591:1584] ,data[1599:1592] ,data[1607:1600] ,data[1799:1792] ,data[1807:1800] ,data[1815:1808] ,data[1823:1816] ,data[1831:1824] ,data[2023:2016] ,data[2031:2024] ,data[2039:2032] ,data[2047:2040] ,data[2055:2048] };
end
199 :begin
 dPIn = {data[1135:1128] ,data[1143:1136] ,data[1151:1144] ,data[1159:1152] ,data[1167:1160] ,data[1359:1352] ,data[1367:1360] ,data[1375:1368] ,data[1383:1376] ,data[1391:1384] ,data[1583:1576] ,data[1591:1584] ,data[1599:1592] ,data[1607:1600] ,data[1615:1608] ,data[1807:1800] ,data[1815:1808] ,data[1823:1816] ,data[1831:1824] ,data[1839:1832] ,data[2031:2024] ,data[2039:2032] ,data[2047:2040] ,data[2055:2048] ,data[2063:2056] };
end
200 :begin
 dPIn = {data[1143:1136] ,data[1151:1144] ,data[1159:1152] ,data[1167:1160] ,data[1175:1168] ,data[1367:1360] ,data[1375:1368] ,data[1383:1376] ,data[1391:1384] ,data[1399:1392] ,data[1591:1584] ,data[1599:1592] ,data[1607:1600] ,data[1615:1608] ,data[1623:1616] ,data[1815:1808] ,data[1823:1816] ,data[1831:1824] ,data[1839:1832] ,data[1847:1840] ,data[2039:2032] ,data[2047:2040] ,data[2055:2048] ,data[2063:2056] ,data[2071:2064] };
end
201 :begin
 dPIn = {data[1151:1144] ,data[1159:1152] ,data[1167:1160] ,data[1175:1168] ,data[1183:1176] ,data[1375:1368] ,data[1383:1376] ,data[1391:1384] ,data[1399:1392] ,data[1407:1400] ,data[1599:1592] ,data[1607:1600] ,data[1615:1608] ,data[1623:1616] ,data[1631:1624] ,data[1823:1816] ,data[1831:1824] ,data[1839:1832] ,data[1847:1840] ,data[1855:1848] ,data[2047:2040] ,data[2055:2048] ,data[2063:2056] ,data[2071:2064] ,data[2079:2072] };
end
202 :begin
 dPIn = {data[1159:1152] ,data[1167:1160] ,data[1175:1168] ,data[1183:1176] ,data[1191:1184] ,data[1383:1376] ,data[1391:1384] ,data[1399:1392] ,data[1407:1400] ,data[1415:1408] ,data[1607:1600] ,data[1615:1608] ,data[1623:1616] ,data[1631:1624] ,data[1639:1632] ,data[1831:1824] ,data[1839:1832] ,data[1847:1840] ,data[1855:1848] ,data[1863:1856] ,data[2055:2048] ,data[2063:2056] ,data[2071:2064] ,data[2079:2072] ,data[2087:2080] };
end
203 :begin
 dPIn = {data[1167:1160] ,data[1175:1168] ,data[1183:1176] ,data[1191:1184] ,data[1199:1192] ,data[1391:1384] ,data[1399:1392] ,data[1407:1400] ,data[1415:1408] ,data[1423:1416] ,data[1615:1608] ,data[1623:1616] ,data[1631:1624] ,data[1639:1632] ,data[1647:1640] ,data[1839:1832] ,data[1847:1840] ,data[1855:1848] ,data[1863:1856] ,data[1871:1864] ,data[2063:2056] ,data[2071:2064] ,data[2079:2072] ,data[2087:2080] ,data[2095:2088] };
end
204 :begin
 dPIn = {data[1175:1168] ,data[1183:1176] ,data[1191:1184] ,data[1199:1192] ,data[1207:1200] ,data[1399:1392] ,data[1407:1400] ,data[1415:1408] ,data[1423:1416] ,data[1431:1424] ,data[1623:1616] ,data[1631:1624] ,data[1639:1632] ,data[1647:1640] ,data[1655:1648] ,data[1847:1840] ,data[1855:1848] ,data[1863:1856] ,data[1871:1864] ,data[1879:1872] ,data[2071:2064] ,data[2079:2072] ,data[2087:2080] ,data[2095:2088] ,data[2103:2096] };
end
205 :begin
 dPIn = {data[1183:1176] ,data[1191:1184] ,data[1199:1192] ,data[1207:1200] ,data[1215:1208] ,data[1407:1400] ,data[1415:1408] ,data[1423:1416] ,data[1431:1424] ,data[1439:1432] ,data[1631:1624] ,data[1639:1632] ,data[1647:1640] ,data[1655:1648] ,data[1663:1656] ,data[1855:1848] ,data[1863:1856] ,data[1871:1864] ,data[1879:1872] ,data[1887:1880] ,data[2079:2072] ,data[2087:2080] ,data[2095:2088] ,data[2103:2096] ,data[2111:2104] };
end
206 :begin
 dPIn = {data[1191:1184] ,data[1199:1192] ,data[1207:1200] ,data[1215:1208] ,data[1223:1216] ,data[1415:1408] ,data[1423:1416] ,data[1431:1424] ,data[1439:1432] ,data[1447:1440] ,data[1639:1632] ,data[1647:1640] ,data[1655:1648] ,data[1663:1656] ,data[1671:1664] ,data[1863:1856] ,data[1871:1864] ,data[1879:1872] ,data[1887:1880] ,data[1895:1888] ,data[2087:2080] ,data[2095:2088] ,data[2103:2096] ,data[2111:2104] ,data[2119:2112] };
end
207 :begin
 dPIn = {data[1199:1192] ,data[1207:1200] ,data[1215:1208] ,data[1223:1216] ,data[1231:1224] ,data[1423:1416] ,data[1431:1424] ,data[1439:1432] ,data[1447:1440] ,data[1455:1448] ,data[1647:1640] ,data[1655:1648] ,data[1663:1656] ,data[1671:1664] ,data[1679:1672] ,data[1871:1864] ,data[1879:1872] ,data[1887:1880] ,data[1895:1888] ,data[1903:1896] ,data[2095:2088] ,data[2103:2096] ,data[2111:2104] ,data[2119:2112] ,data[2127:2120] };
end
208 :begin
 dPIn = {data[1207:1200] ,data[1215:1208] ,data[1223:1216] ,data[1231:1224] ,data[1239:1232] ,data[1431:1424] ,data[1439:1432] ,data[1447:1440] ,data[1455:1448] ,data[1463:1456] ,data[1655:1648] ,data[1663:1656] ,data[1671:1664] ,data[1679:1672] ,data[1687:1680] ,data[1879:1872] ,data[1887:1880] ,data[1895:1888] ,data[1903:1896] ,data[1911:1904] ,data[2103:2096] ,data[2111:2104] ,data[2119:2112] ,data[2127:2120] ,data[2135:2128] };
end
209 :begin
 dPIn = {data[1215:1208] ,data[1223:1216] ,data[1231:1224] ,data[1239:1232] ,data[1247:1240] ,data[1439:1432] ,data[1447:1440] ,data[1455:1448] ,data[1463:1456] ,data[1471:1464] ,data[1663:1656] ,data[1671:1664] ,data[1679:1672] ,data[1687:1680] ,data[1695:1688] ,data[1887:1880] ,data[1895:1888] ,data[1903:1896] ,data[1911:1904] ,data[1919:1912] ,data[2111:2104] ,data[2119:2112] ,data[2127:2120] ,data[2135:2128] ,data[2143:2136] };
end
210 :begin
 dPIn = {data[1223:1216] ,data[1231:1224] ,data[1239:1232] ,data[1247:1240] ,data[1255:1248] ,data[1447:1440] ,data[1455:1448] ,data[1463:1456] ,data[1471:1464] ,data[1479:1472] ,data[1671:1664] ,data[1679:1672] ,data[1687:1680] ,data[1695:1688] ,data[1703:1696] ,data[1895:1888] ,data[1903:1896] ,data[1911:1904] ,data[1919:1912] ,data[1927:1920] ,data[2119:2112] ,data[2127:2120] ,data[2135:2128] ,data[2143:2136] ,data[2151:2144] };
end
211 :begin
 dPIn = {data[1231:1224] ,data[1239:1232] ,data[1247:1240] ,data[1255:1248] ,data[1263:1256] ,data[1455:1448] ,data[1463:1456] ,data[1471:1464] ,data[1479:1472] ,data[1487:1480] ,data[1679:1672] ,data[1687:1680] ,data[1695:1688] ,data[1703:1696] ,data[1711:1704] ,data[1903:1896] ,data[1911:1904] ,data[1919:1912] ,data[1927:1920] ,data[1935:1928] ,data[2127:2120] ,data[2135:2128] ,data[2143:2136] ,data[2151:2144] ,data[2159:2152] };
end
212 :begin
 dPIn = {data[1239:1232] ,data[1247:1240] ,data[1255:1248] ,data[1263:1256] ,data[1271:1264] ,data[1463:1456] ,data[1471:1464] ,data[1479:1472] ,data[1487:1480] ,data[1495:1488] ,data[1687:1680] ,data[1695:1688] ,data[1703:1696] ,data[1711:1704] ,data[1719:1712] ,data[1911:1904] ,data[1919:1912] ,data[1927:1920] ,data[1935:1928] ,data[1943:1936] ,data[2135:2128] ,data[2143:2136] ,data[2151:2144] ,data[2159:2152] ,data[2167:2160] };
end
213 :begin
 dPIn = {data[1247:1240] ,data[1255:1248] ,data[1263:1256] ,data[1271:1264] ,data[1279:1272] ,data[1471:1464] ,data[1479:1472] ,data[1487:1480] ,data[1495:1488] ,data[1503:1496] ,data[1695:1688] ,data[1703:1696] ,data[1711:1704] ,data[1719:1712] ,data[1727:1720] ,data[1919:1912] ,data[1927:1920] ,data[1935:1928] ,data[1943:1936] ,data[1951:1944] ,data[2143:2136] ,data[2151:2144] ,data[2159:2152] ,data[2167:2160] ,data[2175:2168] };
end
214 :begin
 dPIn = {data[1255:1248] ,data[1263:1256] ,data[1271:1264] ,data[1279:1272] ,data[1287:1280] ,data[1479:1472] ,data[1487:1480] ,data[1495:1488] ,data[1503:1496] ,data[1511:1504] ,data[1703:1696] ,data[1711:1704] ,data[1719:1712] ,data[1727:1720] ,data[1735:1728] ,data[1927:1920] ,data[1935:1928] ,data[1943:1936] ,data[1951:1944] ,data[1959:1952] ,data[2151:2144] ,data[2159:2152] ,data[2167:2160] ,data[2175:2168] ,data[2183:2176] };
end
215 :begin
 dPIn = {data[1263:1256] ,data[1271:1264] ,data[1279:1272] ,data[1287:1280] ,data[1295:1288] ,data[1487:1480] ,data[1495:1488] ,data[1503:1496] ,data[1511:1504] ,data[1519:1512] ,data[1711:1704] ,data[1719:1712] ,data[1727:1720] ,data[1735:1728] ,data[1743:1736] ,data[1935:1928] ,data[1943:1936] ,data[1951:1944] ,data[1959:1952] ,data[1967:1960] ,data[2159:2152] ,data[2167:2160] ,data[2175:2168] ,data[2183:2176] ,data[2191:2184] };
end
216 :begin
 dPIn = {data[1271:1264] ,data[1279:1272] ,data[1287:1280] ,data[1295:1288] ,data[1303:1296] ,data[1495:1488] ,data[1503:1496] ,data[1511:1504] ,data[1519:1512] ,data[1527:1520] ,data[1719:1712] ,data[1727:1720] ,data[1735:1728] ,data[1743:1736] ,data[1751:1744] ,data[1943:1936] ,data[1951:1944] ,data[1959:1952] ,data[1967:1960] ,data[1975:1968] ,data[2167:2160] ,data[2175:2168] ,data[2183:2176] ,data[2191:2184] ,data[2199:2192] };
end
217 :begin
 dPIn = {data[1279:1272] ,data[1287:1280] ,data[1295:1288] ,data[1303:1296] ,data[1311:1304] ,data[1503:1496] ,data[1511:1504] ,data[1519:1512] ,data[1527:1520] ,data[1535:1528] ,data[1727:1720] ,data[1735:1728] ,data[1743:1736] ,data[1751:1744] ,data[1759:1752] ,data[1951:1944] ,data[1959:1952] ,data[1967:1960] ,data[1975:1968] ,data[1983:1976] ,data[2175:2168] ,data[2183:2176] ,data[2191:2184] ,data[2199:2192] ,data[2207:2200] };
end
218 :begin
 dPIn = {data[1287:1280] ,data[1295:1288] ,data[1303:1296] ,data[1311:1304] ,data[1319:1312] ,data[1511:1504] ,data[1519:1512] ,data[1527:1520] ,data[1535:1528] ,data[1543:1536] ,data[1735:1728] ,data[1743:1736] ,data[1751:1744] ,data[1759:1752] ,data[1767:1760] ,data[1959:1952] ,data[1967:1960] ,data[1975:1968] ,data[1983:1976] ,data[1991:1984] ,data[2183:2176] ,data[2191:2184] ,data[2199:2192] ,data[2207:2200] ,data[2215:2208] };
end
219 :begin
 dPIn = {data[1295:1288] ,data[1303:1296] ,data[1311:1304] ,data[1319:1312] ,data[1327:1320] ,data[1519:1512] ,data[1527:1520] ,data[1535:1528] ,data[1543:1536] ,data[1551:1544] ,data[1743:1736] ,data[1751:1744] ,data[1759:1752] ,data[1767:1760] ,data[1775:1768] ,data[1967:1960] ,data[1975:1968] ,data[1983:1976] ,data[1991:1984] ,data[1999:1992] ,data[2191:2184] ,data[2199:2192] ,data[2207:2200] ,data[2215:2208] ,data[2223:2216] };
end
220 :begin
 dPIn = {data[1303:1296] ,data[1311:1304] ,data[1319:1312] ,data[1327:1320] ,data[1335:1328] ,data[1527:1520] ,data[1535:1528] ,data[1543:1536] ,data[1551:1544] ,data[1559:1552] ,data[1751:1744] ,data[1759:1752] ,data[1767:1760] ,data[1775:1768] ,data[1783:1776] ,data[1975:1968] ,data[1983:1976] ,data[1991:1984] ,data[1999:1992] ,data[2007:2000] ,data[2199:2192] ,data[2207:2200] ,data[2215:2208] ,data[2223:2216] ,data[2231:2224] };
end
221 :begin
 dPIn = {data[1311:1304] ,data[1319:1312] ,data[1327:1320] ,data[1335:1328] ,data[1343:1336] ,data[1535:1528] ,data[1543:1536] ,data[1551:1544] ,data[1559:1552] ,data[1567:1560] ,data[1759:1752] ,data[1767:1760] ,data[1775:1768] ,data[1783:1776] ,data[1791:1784] ,data[1983:1976] ,data[1991:1984] ,data[1999:1992] ,data[2007:2000] ,data[2015:2008] ,data[2207:2200] ,data[2215:2208] ,data[2223:2216] ,data[2231:2224] ,data[2239:2232] };
end
222 :begin
 dPIn = {data[1319:1312] ,data[1327:1320] ,data[1335:1328] ,data[1343:1336] ,0 ,data[1543:1536] ,data[1551:1544] ,data[1559:1552] ,data[1567:1560] ,0 ,data[1767:1760] ,data[1775:1768] ,data[1783:1776] ,data[1791:1784] ,0 ,data[1991:1984] ,data[1999:1992] ,data[2007:2000] ,data[2015:2008] ,0 ,data[2215:2208] ,data[2223:2216] ,data[2231:2224] ,data[2239:2232] ,0 };
end
223 :begin
 dPIn = {data[1327:1320] ,data[1335:1328] ,data[1343:1336] ,0 ,0 ,data[1551:1544] ,data[1559:1552] ,data[1567:1560] ,0 ,0 ,data[1775:1768] ,data[1783:1776] ,data[1791:1784] ,0 ,0 ,data[1999:1992] ,data[2007:2000] ,data[2015:2008] ,0 ,0 ,data[2223:2216] ,data[2231:2224] ,data[2239:2232] ,0 ,0 };
end
224 :begin
 dPIn = {0 ,0 ,data[1351:1344] ,data[1359:1352] ,data[1367:1360] ,0 ,0 ,data[1575:1568] ,data[1583:1576] ,data[1591:1584] ,0 ,0 ,data[1799:1792] ,data[1807:1800] ,data[1815:1808] ,0 ,0 ,data[2023:2016] ,data[2031:2024] ,data[2039:2032] ,0 ,0 ,data[2247:2240] ,data[2255:2248] ,data[2263:2256] };
end
225 :begin
 dPIn = {0 ,data[1351:1344] ,data[1359:1352] ,data[1367:1360] ,data[1375:1368] ,0 ,data[1575:1568] ,data[1583:1576] ,data[1591:1584] ,data[1599:1592] ,0 ,data[1799:1792] ,data[1807:1800] ,data[1815:1808] ,data[1823:1816] ,0 ,data[2023:2016] ,data[2031:2024] ,data[2039:2032] ,data[2047:2040] ,0 ,data[2247:2240] ,data[2255:2248] ,data[2263:2256] ,data[2271:2264] };
end
226 :begin
 dPIn = {data[1351:1344] ,data[1359:1352] ,data[1367:1360] ,data[1375:1368] ,data[1383:1376] ,data[1575:1568] ,data[1583:1576] ,data[1591:1584] ,data[1599:1592] ,data[1607:1600] ,data[1799:1792] ,data[1807:1800] ,data[1815:1808] ,data[1823:1816] ,data[1831:1824] ,data[2023:2016] ,data[2031:2024] ,data[2039:2032] ,data[2047:2040] ,data[2055:2048] ,data[2247:2240] ,data[2255:2248] ,data[2263:2256] ,data[2271:2264] ,data[2279:2272] };
end
227 :begin
 dPIn = {data[1359:1352] ,data[1367:1360] ,data[1375:1368] ,data[1383:1376] ,data[1391:1384] ,data[1583:1576] ,data[1591:1584] ,data[1599:1592] ,data[1607:1600] ,data[1615:1608] ,data[1807:1800] ,data[1815:1808] ,data[1823:1816] ,data[1831:1824] ,data[1839:1832] ,data[2031:2024] ,data[2039:2032] ,data[2047:2040] ,data[2055:2048] ,data[2063:2056] ,data[2255:2248] ,data[2263:2256] ,data[2271:2264] ,data[2279:2272] ,data[2287:2280] };
end
228 :begin
 dPIn = {data[1367:1360] ,data[1375:1368] ,data[1383:1376] ,data[1391:1384] ,data[1399:1392] ,data[1591:1584] ,data[1599:1592] ,data[1607:1600] ,data[1615:1608] ,data[1623:1616] ,data[1815:1808] ,data[1823:1816] ,data[1831:1824] ,data[1839:1832] ,data[1847:1840] ,data[2039:2032] ,data[2047:2040] ,data[2055:2048] ,data[2063:2056] ,data[2071:2064] ,data[2263:2256] ,data[2271:2264] ,data[2279:2272] ,data[2287:2280] ,data[2295:2288] };
end
229 :begin
 dPIn = {data[1375:1368] ,data[1383:1376] ,data[1391:1384] ,data[1399:1392] ,data[1407:1400] ,data[1599:1592] ,data[1607:1600] ,data[1615:1608] ,data[1623:1616] ,data[1631:1624] ,data[1823:1816] ,data[1831:1824] ,data[1839:1832] ,data[1847:1840] ,data[1855:1848] ,data[2047:2040] ,data[2055:2048] ,data[2063:2056] ,data[2071:2064] ,data[2079:2072] ,data[2271:2264] ,data[2279:2272] ,data[2287:2280] ,data[2295:2288] ,data[2303:2296] };
end
230 :begin
 dPIn = {data[1383:1376] ,data[1391:1384] ,data[1399:1392] ,data[1407:1400] ,data[1415:1408] ,data[1607:1600] ,data[1615:1608] ,data[1623:1616] ,data[1631:1624] ,data[1639:1632] ,data[1831:1824] ,data[1839:1832] ,data[1847:1840] ,data[1855:1848] ,data[1863:1856] ,data[2055:2048] ,data[2063:2056] ,data[2071:2064] ,data[2079:2072] ,data[2087:2080] ,data[2279:2272] ,data[2287:2280] ,data[2295:2288] ,data[2303:2296] ,data[2311:2304] };
end
231 :begin
 dPIn = {data[1391:1384] ,data[1399:1392] ,data[1407:1400] ,data[1415:1408] ,data[1423:1416] ,data[1615:1608] ,data[1623:1616] ,data[1631:1624] ,data[1639:1632] ,data[1647:1640] ,data[1839:1832] ,data[1847:1840] ,data[1855:1848] ,data[1863:1856] ,data[1871:1864] ,data[2063:2056] ,data[2071:2064] ,data[2079:2072] ,data[2087:2080] ,data[2095:2088] ,data[2287:2280] ,data[2295:2288] ,data[2303:2296] ,data[2311:2304] ,data[2319:2312] };
end
232 :begin
 dPIn = {data[1399:1392] ,data[1407:1400] ,data[1415:1408] ,data[1423:1416] ,data[1431:1424] ,data[1623:1616] ,data[1631:1624] ,data[1639:1632] ,data[1647:1640] ,data[1655:1648] ,data[1847:1840] ,data[1855:1848] ,data[1863:1856] ,data[1871:1864] ,data[1879:1872] ,data[2071:2064] ,data[2079:2072] ,data[2087:2080] ,data[2095:2088] ,data[2103:2096] ,data[2295:2288] ,data[2303:2296] ,data[2311:2304] ,data[2319:2312] ,data[2327:2320] };
end
233 :begin
 dPIn = {data[1407:1400] ,data[1415:1408] ,data[1423:1416] ,data[1431:1424] ,data[1439:1432] ,data[1631:1624] ,data[1639:1632] ,data[1647:1640] ,data[1655:1648] ,data[1663:1656] ,data[1855:1848] ,data[1863:1856] ,data[1871:1864] ,data[1879:1872] ,data[1887:1880] ,data[2079:2072] ,data[2087:2080] ,data[2095:2088] ,data[2103:2096] ,data[2111:2104] ,data[2303:2296] ,data[2311:2304] ,data[2319:2312] ,data[2327:2320] ,data[2335:2328] };
end
234 :begin
 dPIn = {data[1415:1408] ,data[1423:1416] ,data[1431:1424] ,data[1439:1432] ,data[1447:1440] ,data[1639:1632] ,data[1647:1640] ,data[1655:1648] ,data[1663:1656] ,data[1671:1664] ,data[1863:1856] ,data[1871:1864] ,data[1879:1872] ,data[1887:1880] ,data[1895:1888] ,data[2087:2080] ,data[2095:2088] ,data[2103:2096] ,data[2111:2104] ,data[2119:2112] ,data[2311:2304] ,data[2319:2312] ,data[2327:2320] ,data[2335:2328] ,data[2343:2336] };
end
235 :begin
 dPIn = {data[1423:1416] ,data[1431:1424] ,data[1439:1432] ,data[1447:1440] ,data[1455:1448] ,data[1647:1640] ,data[1655:1648] ,data[1663:1656] ,data[1671:1664] ,data[1679:1672] ,data[1871:1864] ,data[1879:1872] ,data[1887:1880] ,data[1895:1888] ,data[1903:1896] ,data[2095:2088] ,data[2103:2096] ,data[2111:2104] ,data[2119:2112] ,data[2127:2120] ,data[2319:2312] ,data[2327:2320] ,data[2335:2328] ,data[2343:2336] ,data[2351:2344] };
end
236 :begin
 dPIn = {data[1431:1424] ,data[1439:1432] ,data[1447:1440] ,data[1455:1448] ,data[1463:1456] ,data[1655:1648] ,data[1663:1656] ,data[1671:1664] ,data[1679:1672] ,data[1687:1680] ,data[1879:1872] ,data[1887:1880] ,data[1895:1888] ,data[1903:1896] ,data[1911:1904] ,data[2103:2096] ,data[2111:2104] ,data[2119:2112] ,data[2127:2120] ,data[2135:2128] ,data[2327:2320] ,data[2335:2328] ,data[2343:2336] ,data[2351:2344] ,data[2359:2352] };
end
237 :begin
 dPIn = {data[1439:1432] ,data[1447:1440] ,data[1455:1448] ,data[1463:1456] ,data[1471:1464] ,data[1663:1656] ,data[1671:1664] ,data[1679:1672] ,data[1687:1680] ,data[1695:1688] ,data[1887:1880] ,data[1895:1888] ,data[1903:1896] ,data[1911:1904] ,data[1919:1912] ,data[2111:2104] ,data[2119:2112] ,data[2127:2120] ,data[2135:2128] ,data[2143:2136] ,data[2335:2328] ,data[2343:2336] ,data[2351:2344] ,data[2359:2352] ,data[2367:2360] };
end
238 :begin
 dPIn = {data[1447:1440] ,data[1455:1448] ,data[1463:1456] ,data[1471:1464] ,data[1479:1472] ,data[1671:1664] ,data[1679:1672] ,data[1687:1680] ,data[1695:1688] ,data[1703:1696] ,data[1895:1888] ,data[1903:1896] ,data[1911:1904] ,data[1919:1912] ,data[1927:1920] ,data[2119:2112] ,data[2127:2120] ,data[2135:2128] ,data[2143:2136] ,data[2151:2144] ,data[2343:2336] ,data[2351:2344] ,data[2359:2352] ,data[2367:2360] ,data[2375:2368] };
end
239 :begin
 dPIn = {data[1455:1448] ,data[1463:1456] ,data[1471:1464] ,data[1479:1472] ,data[1487:1480] ,data[1679:1672] ,data[1687:1680] ,data[1695:1688] ,data[1703:1696] ,data[1711:1704] ,data[1903:1896] ,data[1911:1904] ,data[1919:1912] ,data[1927:1920] ,data[1935:1928] ,data[2127:2120] ,data[2135:2128] ,data[2143:2136] ,data[2151:2144] ,data[2159:2152] ,data[2351:2344] ,data[2359:2352] ,data[2367:2360] ,data[2375:2368] ,data[2383:2376] };
end
240 :begin
 dPIn = {data[1463:1456] ,data[1471:1464] ,data[1479:1472] ,data[1487:1480] ,data[1495:1488] ,data[1687:1680] ,data[1695:1688] ,data[1703:1696] ,data[1711:1704] ,data[1719:1712] ,data[1911:1904] ,data[1919:1912] ,data[1927:1920] ,data[1935:1928] ,data[1943:1936] ,data[2135:2128] ,data[2143:2136] ,data[2151:2144] ,data[2159:2152] ,data[2167:2160] ,data[2359:2352] ,data[2367:2360] ,data[2375:2368] ,data[2383:2376] ,data[2391:2384] };
end
241 :begin
 dPIn = {data[1471:1464] ,data[1479:1472] ,data[1487:1480] ,data[1495:1488] ,data[1503:1496] ,data[1695:1688] ,data[1703:1696] ,data[1711:1704] ,data[1719:1712] ,data[1727:1720] ,data[1919:1912] ,data[1927:1920] ,data[1935:1928] ,data[1943:1936] ,data[1951:1944] ,data[2143:2136] ,data[2151:2144] ,data[2159:2152] ,data[2167:2160] ,data[2175:2168] ,data[2367:2360] ,data[2375:2368] ,data[2383:2376] ,data[2391:2384] ,data[2399:2392] };
end
242 :begin
 dPIn = {data[1479:1472] ,data[1487:1480] ,data[1495:1488] ,data[1503:1496] ,data[1511:1504] ,data[1703:1696] ,data[1711:1704] ,data[1719:1712] ,data[1727:1720] ,data[1735:1728] ,data[1927:1920] ,data[1935:1928] ,data[1943:1936] ,data[1951:1944] ,data[1959:1952] ,data[2151:2144] ,data[2159:2152] ,data[2167:2160] ,data[2175:2168] ,data[2183:2176] ,data[2375:2368] ,data[2383:2376] ,data[2391:2384] ,data[2399:2392] ,data[2407:2400] };
end
243 :begin
 dPIn = {data[1487:1480] ,data[1495:1488] ,data[1503:1496] ,data[1511:1504] ,data[1519:1512] ,data[1711:1704] ,data[1719:1712] ,data[1727:1720] ,data[1735:1728] ,data[1743:1736] ,data[1935:1928] ,data[1943:1936] ,data[1951:1944] ,data[1959:1952] ,data[1967:1960] ,data[2159:2152] ,data[2167:2160] ,data[2175:2168] ,data[2183:2176] ,data[2191:2184] ,data[2383:2376] ,data[2391:2384] ,data[2399:2392] ,data[2407:2400] ,data[2415:2408] };
end
244 :begin
 dPIn = {data[1495:1488] ,data[1503:1496] ,data[1511:1504] ,data[1519:1512] ,data[1527:1520] ,data[1719:1712] ,data[1727:1720] ,data[1735:1728] ,data[1743:1736] ,data[1751:1744] ,data[1943:1936] ,data[1951:1944] ,data[1959:1952] ,data[1967:1960] ,data[1975:1968] ,data[2167:2160] ,data[2175:2168] ,data[2183:2176] ,data[2191:2184] ,data[2199:2192] ,data[2391:2384] ,data[2399:2392] ,data[2407:2400] ,data[2415:2408] ,data[2423:2416] };
end
245 :begin
 dPIn = {data[1503:1496] ,data[1511:1504] ,data[1519:1512] ,data[1527:1520] ,data[1535:1528] ,data[1727:1720] ,data[1735:1728] ,data[1743:1736] ,data[1751:1744] ,data[1759:1752] ,data[1951:1944] ,data[1959:1952] ,data[1967:1960] ,data[1975:1968] ,data[1983:1976] ,data[2175:2168] ,data[2183:2176] ,data[2191:2184] ,data[2199:2192] ,data[2207:2200] ,data[2399:2392] ,data[2407:2400] ,data[2415:2408] ,data[2423:2416] ,data[2431:2424] };
end
246 :begin
 dPIn = {data[1511:1504] ,data[1519:1512] ,data[1527:1520] ,data[1535:1528] ,data[1543:1536] ,data[1735:1728] ,data[1743:1736] ,data[1751:1744] ,data[1759:1752] ,data[1767:1760] ,data[1959:1952] ,data[1967:1960] ,data[1975:1968] ,data[1983:1976] ,data[1991:1984] ,data[2183:2176] ,data[2191:2184] ,data[2199:2192] ,data[2207:2200] ,data[2215:2208] ,data[2407:2400] ,data[2415:2408] ,data[2423:2416] ,data[2431:2424] ,data[2439:2432] };
end
247 :begin
 dPIn = {data[1519:1512] ,data[1527:1520] ,data[1535:1528] ,data[1543:1536] ,data[1551:1544] ,data[1743:1736] ,data[1751:1744] ,data[1759:1752] ,data[1767:1760] ,data[1775:1768] ,data[1967:1960] ,data[1975:1968] ,data[1983:1976] ,data[1991:1984] ,data[1999:1992] ,data[2191:2184] ,data[2199:2192] ,data[2207:2200] ,data[2215:2208] ,data[2223:2216] ,data[2415:2408] ,data[2423:2416] ,data[2431:2424] ,data[2439:2432] ,data[2447:2440] };
end
248 :begin
 dPIn = {data[1527:1520] ,data[1535:1528] ,data[1543:1536] ,data[1551:1544] ,data[1559:1552] ,data[1751:1744] ,data[1759:1752] ,data[1767:1760] ,data[1775:1768] ,data[1783:1776] ,data[1975:1968] ,data[1983:1976] ,data[1991:1984] ,data[1999:1992] ,data[2007:2000] ,data[2199:2192] ,data[2207:2200] ,data[2215:2208] ,data[2223:2216] ,data[2231:2224] ,data[2423:2416] ,data[2431:2424] ,data[2439:2432] ,data[2447:2440] ,data[2455:2448] };
end
249 :begin
 dPIn = {data[1535:1528] ,data[1543:1536] ,data[1551:1544] ,data[1559:1552] ,data[1567:1560] ,data[1759:1752] ,data[1767:1760] ,data[1775:1768] ,data[1783:1776] ,data[1791:1784] ,data[1983:1976] ,data[1991:1984] ,data[1999:1992] ,data[2007:2000] ,data[2015:2008] ,data[2207:2200] ,data[2215:2208] ,data[2223:2216] ,data[2231:2224] ,data[2239:2232] ,data[2431:2424] ,data[2439:2432] ,data[2447:2440] ,data[2455:2448] ,data[2463:2456] };
end
250 :begin
 dPIn = {data[1543:1536] ,data[1551:1544] ,data[1559:1552] ,data[1567:1560] ,0 ,data[1767:1760] ,data[1775:1768] ,data[1783:1776] ,data[1791:1784] ,0 ,data[1991:1984] ,data[1999:1992] ,data[2007:2000] ,data[2015:2008] ,0 ,data[2215:2208] ,data[2223:2216] ,data[2231:2224] ,data[2239:2232] ,0 ,data[2439:2432] ,data[2447:2440] ,data[2455:2448] ,data[2463:2456] ,0 };
end
251 :begin
 dPIn = {data[1551:1544] ,data[1559:1552] ,data[1567:1560] ,0 ,0 ,data[1775:1768] ,data[1783:1776] ,data[1791:1784] ,0 ,0 ,data[1999:1992] ,data[2007:2000] ,data[2015:2008] ,0 ,0 ,data[2223:2216] ,data[2231:2224] ,data[2239:2232] ,0 ,0 ,data[2447:2440] ,data[2455:2448] ,data[2463:2456] ,0 ,0 };
end
252 :begin
 dPIn = {0 ,0 ,data[1575:1568] ,data[1583:1576] ,data[1591:1584] ,0 ,0 ,data[1799:1792] ,data[1807:1800] ,data[1815:1808] ,0 ,0 ,data[2023:2016] ,data[2031:2024] ,data[2039:2032] ,0 ,0 ,data[2247:2240] ,data[2255:2248] ,data[2263:2256] ,0 ,0 ,data[2471:2464] ,data[2479:2472] ,data[2487:2480] };
end
253 :begin
 dPIn = {0 ,data[1575:1568] ,data[1583:1576] ,data[1591:1584] ,data[1599:1592] ,0 ,data[1799:1792] ,data[1807:1800] ,data[1815:1808] ,data[1823:1816] ,0 ,data[2023:2016] ,data[2031:2024] ,data[2039:2032] ,data[2047:2040] ,0 ,data[2247:2240] ,data[2255:2248] ,data[2263:2256] ,data[2271:2264] ,0 ,data[2471:2464] ,data[2479:2472] ,data[2487:2480] ,data[2495:2488] };
end
254 :begin
 dPIn = {data[1575:1568] ,data[1583:1576] ,data[1591:1584] ,data[1599:1592] ,data[1607:1600] ,data[1799:1792] ,data[1807:1800] ,data[1815:1808] ,data[1823:1816] ,data[1831:1824] ,data[2023:2016] ,data[2031:2024] ,data[2039:2032] ,data[2047:2040] ,data[2055:2048] ,data[2247:2240] ,data[2255:2248] ,data[2263:2256] ,data[2271:2264] ,data[2279:2272] ,data[2471:2464] ,data[2479:2472] ,data[2487:2480] ,data[2495:2488] ,data[2503:2496] };
end
255 :begin
 dPIn = {data[1583:1576] ,data[1591:1584] ,data[1599:1592] ,data[1607:1600] ,data[1615:1608] ,data[1807:1800] ,data[1815:1808] ,data[1823:1816] ,data[1831:1824] ,data[1839:1832] ,data[2031:2024] ,data[2039:2032] ,data[2047:2040] ,data[2055:2048] ,data[2063:2056] ,data[2255:2248] ,data[2263:2256] ,data[2271:2264] ,data[2279:2272] ,data[2287:2280] ,data[2479:2472] ,data[2487:2480] ,data[2495:2488] ,data[2503:2496] ,data[2511:2504] };
end
256 :begin
 dPIn = {data[1591:1584] ,data[1599:1592] ,data[1607:1600] ,data[1615:1608] ,data[1623:1616] ,data[1815:1808] ,data[1823:1816] ,data[1831:1824] ,data[1839:1832] ,data[1847:1840] ,data[2039:2032] ,data[2047:2040] ,data[2055:2048] ,data[2063:2056] ,data[2071:2064] ,data[2263:2256] ,data[2271:2264] ,data[2279:2272] ,data[2287:2280] ,data[2295:2288] ,data[2487:2480] ,data[2495:2488] ,data[2503:2496] ,data[2511:2504] ,data[2519:2512] };
end
257 :begin
 dPIn = {data[1599:1592] ,data[1607:1600] ,data[1615:1608] ,data[1623:1616] ,data[1631:1624] ,data[1823:1816] ,data[1831:1824] ,data[1839:1832] ,data[1847:1840] ,data[1855:1848] ,data[2047:2040] ,data[2055:2048] ,data[2063:2056] ,data[2071:2064] ,data[2079:2072] ,data[2271:2264] ,data[2279:2272] ,data[2287:2280] ,data[2295:2288] ,data[2303:2296] ,data[2495:2488] ,data[2503:2496] ,data[2511:2504] ,data[2519:2512] ,data[2527:2520] };
end
258 :begin
 dPIn = {data[1607:1600] ,data[1615:1608] ,data[1623:1616] ,data[1631:1624] ,data[1639:1632] ,data[1831:1824] ,data[1839:1832] ,data[1847:1840] ,data[1855:1848] ,data[1863:1856] ,data[2055:2048] ,data[2063:2056] ,data[2071:2064] ,data[2079:2072] ,data[2087:2080] ,data[2279:2272] ,data[2287:2280] ,data[2295:2288] ,data[2303:2296] ,data[2311:2304] ,data[2503:2496] ,data[2511:2504] ,data[2519:2512] ,data[2527:2520] ,data[2535:2528] };
end
259 :begin
 dPIn = {data[1615:1608] ,data[1623:1616] ,data[1631:1624] ,data[1639:1632] ,data[1647:1640] ,data[1839:1832] ,data[1847:1840] ,data[1855:1848] ,data[1863:1856] ,data[1871:1864] ,data[2063:2056] ,data[2071:2064] ,data[2079:2072] ,data[2087:2080] ,data[2095:2088] ,data[2287:2280] ,data[2295:2288] ,data[2303:2296] ,data[2311:2304] ,data[2319:2312] ,data[2511:2504] ,data[2519:2512] ,data[2527:2520] ,data[2535:2528] ,data[2543:2536] };
end
260 :begin
 dPIn = {data[1623:1616] ,data[1631:1624] ,data[1639:1632] ,data[1647:1640] ,data[1655:1648] ,data[1847:1840] ,data[1855:1848] ,data[1863:1856] ,data[1871:1864] ,data[1879:1872] ,data[2071:2064] ,data[2079:2072] ,data[2087:2080] ,data[2095:2088] ,data[2103:2096] ,data[2295:2288] ,data[2303:2296] ,data[2311:2304] ,data[2319:2312] ,data[2327:2320] ,data[2519:2512] ,data[2527:2520] ,data[2535:2528] ,data[2543:2536] ,data[2551:2544] };
end
261 :begin
 dPIn = {data[1631:1624] ,data[1639:1632] ,data[1647:1640] ,data[1655:1648] ,data[1663:1656] ,data[1855:1848] ,data[1863:1856] ,data[1871:1864] ,data[1879:1872] ,data[1887:1880] ,data[2079:2072] ,data[2087:2080] ,data[2095:2088] ,data[2103:2096] ,data[2111:2104] ,data[2303:2296] ,data[2311:2304] ,data[2319:2312] ,data[2327:2320] ,data[2335:2328] ,data[2527:2520] ,data[2535:2528] ,data[2543:2536] ,data[2551:2544] ,data[2559:2552] };
end
262 :begin
 dPIn = {data[1639:1632] ,data[1647:1640] ,data[1655:1648] ,data[1663:1656] ,data[1671:1664] ,data[1863:1856] ,data[1871:1864] ,data[1879:1872] ,data[1887:1880] ,data[1895:1888] ,data[2087:2080] ,data[2095:2088] ,data[2103:2096] ,data[2111:2104] ,data[2119:2112] ,data[2311:2304] ,data[2319:2312] ,data[2327:2320] ,data[2335:2328] ,data[2343:2336] ,data[2535:2528] ,data[2543:2536] ,data[2551:2544] ,data[2559:2552] ,data[2567:2560] };
end
263 :begin
 dPIn = {data[1647:1640] ,data[1655:1648] ,data[1663:1656] ,data[1671:1664] ,data[1679:1672] ,data[1871:1864] ,data[1879:1872] ,data[1887:1880] ,data[1895:1888] ,data[1903:1896] ,data[2095:2088] ,data[2103:2096] ,data[2111:2104] ,data[2119:2112] ,data[2127:2120] ,data[2319:2312] ,data[2327:2320] ,data[2335:2328] ,data[2343:2336] ,data[2351:2344] ,data[2543:2536] ,data[2551:2544] ,data[2559:2552] ,data[2567:2560] ,data[2575:2568] };
end
264 :begin
 dPIn = {data[1655:1648] ,data[1663:1656] ,data[1671:1664] ,data[1679:1672] ,data[1687:1680] ,data[1879:1872] ,data[1887:1880] ,data[1895:1888] ,data[1903:1896] ,data[1911:1904] ,data[2103:2096] ,data[2111:2104] ,data[2119:2112] ,data[2127:2120] ,data[2135:2128] ,data[2327:2320] ,data[2335:2328] ,data[2343:2336] ,data[2351:2344] ,data[2359:2352] ,data[2551:2544] ,data[2559:2552] ,data[2567:2560] ,data[2575:2568] ,data[2583:2576] };
end
265 :begin
 dPIn = {data[1663:1656] ,data[1671:1664] ,data[1679:1672] ,data[1687:1680] ,data[1695:1688] ,data[1887:1880] ,data[1895:1888] ,data[1903:1896] ,data[1911:1904] ,data[1919:1912] ,data[2111:2104] ,data[2119:2112] ,data[2127:2120] ,data[2135:2128] ,data[2143:2136] ,data[2335:2328] ,data[2343:2336] ,data[2351:2344] ,data[2359:2352] ,data[2367:2360] ,data[2559:2552] ,data[2567:2560] ,data[2575:2568] ,data[2583:2576] ,data[2591:2584] };
end
266 :begin
 dPIn = {data[1671:1664] ,data[1679:1672] ,data[1687:1680] ,data[1695:1688] ,data[1703:1696] ,data[1895:1888] ,data[1903:1896] ,data[1911:1904] ,data[1919:1912] ,data[1927:1920] ,data[2119:2112] ,data[2127:2120] ,data[2135:2128] ,data[2143:2136] ,data[2151:2144] ,data[2343:2336] ,data[2351:2344] ,data[2359:2352] ,data[2367:2360] ,data[2375:2368] ,data[2567:2560] ,data[2575:2568] ,data[2583:2576] ,data[2591:2584] ,data[2599:2592] };
end
267 :begin
 dPIn = {data[1679:1672] ,data[1687:1680] ,data[1695:1688] ,data[1703:1696] ,data[1711:1704] ,data[1903:1896] ,data[1911:1904] ,data[1919:1912] ,data[1927:1920] ,data[1935:1928] ,data[2127:2120] ,data[2135:2128] ,data[2143:2136] ,data[2151:2144] ,data[2159:2152] ,data[2351:2344] ,data[2359:2352] ,data[2367:2360] ,data[2375:2368] ,data[2383:2376] ,data[2575:2568] ,data[2583:2576] ,data[2591:2584] ,data[2599:2592] ,data[2607:2600] };
end
268 :begin
 dPIn = {data[1687:1680] ,data[1695:1688] ,data[1703:1696] ,data[1711:1704] ,data[1719:1712] ,data[1911:1904] ,data[1919:1912] ,data[1927:1920] ,data[1935:1928] ,data[1943:1936] ,data[2135:2128] ,data[2143:2136] ,data[2151:2144] ,data[2159:2152] ,data[2167:2160] ,data[2359:2352] ,data[2367:2360] ,data[2375:2368] ,data[2383:2376] ,data[2391:2384] ,data[2583:2576] ,data[2591:2584] ,data[2599:2592] ,data[2607:2600] ,data[2615:2608] };
end
269 :begin
 dPIn = {data[1695:1688] ,data[1703:1696] ,data[1711:1704] ,data[1719:1712] ,data[1727:1720] ,data[1919:1912] ,data[1927:1920] ,data[1935:1928] ,data[1943:1936] ,data[1951:1944] ,data[2143:2136] ,data[2151:2144] ,data[2159:2152] ,data[2167:2160] ,data[2175:2168] ,data[2367:2360] ,data[2375:2368] ,data[2383:2376] ,data[2391:2384] ,data[2399:2392] ,data[2591:2584] ,data[2599:2592] ,data[2607:2600] ,data[2615:2608] ,data[2623:2616] };
end
270 :begin
 dPIn = {data[1703:1696] ,data[1711:1704] ,data[1719:1712] ,data[1727:1720] ,data[1735:1728] ,data[1927:1920] ,data[1935:1928] ,data[1943:1936] ,data[1951:1944] ,data[1959:1952] ,data[2151:2144] ,data[2159:2152] ,data[2167:2160] ,data[2175:2168] ,data[2183:2176] ,data[2375:2368] ,data[2383:2376] ,data[2391:2384] ,data[2399:2392] ,data[2407:2400] ,data[2599:2592] ,data[2607:2600] ,data[2615:2608] ,data[2623:2616] ,data[2631:2624] };
end
271 :begin
 dPIn = {data[1711:1704] ,data[1719:1712] ,data[1727:1720] ,data[1735:1728] ,data[1743:1736] ,data[1935:1928] ,data[1943:1936] ,data[1951:1944] ,data[1959:1952] ,data[1967:1960] ,data[2159:2152] ,data[2167:2160] ,data[2175:2168] ,data[2183:2176] ,data[2191:2184] ,data[2383:2376] ,data[2391:2384] ,data[2399:2392] ,data[2407:2400] ,data[2415:2408] ,data[2607:2600] ,data[2615:2608] ,data[2623:2616] ,data[2631:2624] ,data[2639:2632] };
end
272 :begin
 dPIn = {data[1719:1712] ,data[1727:1720] ,data[1735:1728] ,data[1743:1736] ,data[1751:1744] ,data[1943:1936] ,data[1951:1944] ,data[1959:1952] ,data[1967:1960] ,data[1975:1968] ,data[2167:2160] ,data[2175:2168] ,data[2183:2176] ,data[2191:2184] ,data[2199:2192] ,data[2391:2384] ,data[2399:2392] ,data[2407:2400] ,data[2415:2408] ,data[2423:2416] ,data[2615:2608] ,data[2623:2616] ,data[2631:2624] ,data[2639:2632] ,data[2647:2640] };
end
273 :begin
 dPIn = {data[1727:1720] ,data[1735:1728] ,data[1743:1736] ,data[1751:1744] ,data[1759:1752] ,data[1951:1944] ,data[1959:1952] ,data[1967:1960] ,data[1975:1968] ,data[1983:1976] ,data[2175:2168] ,data[2183:2176] ,data[2191:2184] ,data[2199:2192] ,data[2207:2200] ,data[2399:2392] ,data[2407:2400] ,data[2415:2408] ,data[2423:2416] ,data[2431:2424] ,data[2623:2616] ,data[2631:2624] ,data[2639:2632] ,data[2647:2640] ,data[2655:2648] };
end
274 :begin
 dPIn = {data[1735:1728] ,data[1743:1736] ,data[1751:1744] ,data[1759:1752] ,data[1767:1760] ,data[1959:1952] ,data[1967:1960] ,data[1975:1968] ,data[1983:1976] ,data[1991:1984] ,data[2183:2176] ,data[2191:2184] ,data[2199:2192] ,data[2207:2200] ,data[2215:2208] ,data[2407:2400] ,data[2415:2408] ,data[2423:2416] ,data[2431:2424] ,data[2439:2432] ,data[2631:2624] ,data[2639:2632] ,data[2647:2640] ,data[2655:2648] ,data[2663:2656] };
end
275 :begin
 dPIn = {data[1743:1736] ,data[1751:1744] ,data[1759:1752] ,data[1767:1760] ,data[1775:1768] ,data[1967:1960] ,data[1975:1968] ,data[1983:1976] ,data[1991:1984] ,data[1999:1992] ,data[2191:2184] ,data[2199:2192] ,data[2207:2200] ,data[2215:2208] ,data[2223:2216] ,data[2415:2408] ,data[2423:2416] ,data[2431:2424] ,data[2439:2432] ,data[2447:2440] ,data[2639:2632] ,data[2647:2640] ,data[2655:2648] ,data[2663:2656] ,data[2671:2664] };
end
276 :begin
 dPIn = {data[1751:1744] ,data[1759:1752] ,data[1767:1760] ,data[1775:1768] ,data[1783:1776] ,data[1975:1968] ,data[1983:1976] ,data[1991:1984] ,data[1999:1992] ,data[2007:2000] ,data[2199:2192] ,data[2207:2200] ,data[2215:2208] ,data[2223:2216] ,data[2231:2224] ,data[2423:2416] ,data[2431:2424] ,data[2439:2432] ,data[2447:2440] ,data[2455:2448] ,data[2647:2640] ,data[2655:2648] ,data[2663:2656] ,data[2671:2664] ,data[2679:2672] };
end
277 :begin
 dPIn = {data[1759:1752] ,data[1767:1760] ,data[1775:1768] ,data[1783:1776] ,data[1791:1784] ,data[1983:1976] ,data[1991:1984] ,data[1999:1992] ,data[2007:2000] ,data[2015:2008] ,data[2207:2200] ,data[2215:2208] ,data[2223:2216] ,data[2231:2224] ,data[2239:2232] ,data[2431:2424] ,data[2439:2432] ,data[2447:2440] ,data[2455:2448] ,data[2463:2456] ,data[2655:2648] ,data[2663:2656] ,data[2671:2664] ,data[2679:2672] ,data[2687:2680] };
end
278 :begin
 dPIn = {data[1767:1760] ,data[1775:1768] ,data[1783:1776] ,data[1791:1784] ,0 ,data[1991:1984] ,data[1999:1992] ,data[2007:2000] ,data[2015:2008] ,0 ,data[2215:2208] ,data[2223:2216] ,data[2231:2224] ,data[2239:2232] ,0 ,data[2439:2432] ,data[2447:2440] ,data[2455:2448] ,data[2463:2456] ,0 ,data[2663:2656] ,data[2671:2664] ,data[2679:2672] ,data[2687:2680] ,0 };
end
279 :begin
 dPIn = {data[1775:1768] ,data[1783:1776] ,data[1791:1784] ,0 ,0 ,data[1999:1992] ,data[2007:2000] ,data[2015:2008] ,0 ,0 ,data[2223:2216] ,data[2231:2224] ,data[2239:2232] ,0 ,0 ,data[2447:2440] ,data[2455:2448] ,data[2463:2456] ,0 ,0 ,data[2671:2664] ,data[2679:2672] ,data[2687:2680] ,0 ,0 };
end
280 :begin
 dPIn = {0 ,0 ,data[1799:1792] ,data[1807:1800] ,data[1815:1808] ,0 ,0 ,data[2023:2016] ,data[2031:2024] ,data[2039:2032] ,0 ,0 ,data[2247:2240] ,data[2255:2248] ,data[2263:2256] ,0 ,0 ,data[2471:2464] ,data[2479:2472] ,data[2487:2480] ,0 ,0 ,data[2695:2688] ,data[2703:2696] ,data[2711:2704] };
end
281 :begin
 dPIn = {0 ,data[1799:1792] ,data[1807:1800] ,data[1815:1808] ,data[1823:1816] ,0 ,data[2023:2016] ,data[2031:2024] ,data[2039:2032] ,data[2047:2040] ,0 ,data[2247:2240] ,data[2255:2248] ,data[2263:2256] ,data[2271:2264] ,0 ,data[2471:2464] ,data[2479:2472] ,data[2487:2480] ,data[2495:2488] ,0 ,data[2695:2688] ,data[2703:2696] ,data[2711:2704] ,data[2719:2712] };
end
282 :begin
 dPIn = {data[1799:1792] ,data[1807:1800] ,data[1815:1808] ,data[1823:1816] ,data[1831:1824] ,data[2023:2016] ,data[2031:2024] ,data[2039:2032] ,data[2047:2040] ,data[2055:2048] ,data[2247:2240] ,data[2255:2248] ,data[2263:2256] ,data[2271:2264] ,data[2279:2272] ,data[2471:2464] ,data[2479:2472] ,data[2487:2480] ,data[2495:2488] ,data[2503:2496] ,data[2695:2688] ,data[2703:2696] ,data[2711:2704] ,data[2719:2712] ,data[2727:2720] };
end
283 :begin
 dPIn = {data[1807:1800] ,data[1815:1808] ,data[1823:1816] ,data[1831:1824] ,data[1839:1832] ,data[2031:2024] ,data[2039:2032] ,data[2047:2040] ,data[2055:2048] ,data[2063:2056] ,data[2255:2248] ,data[2263:2256] ,data[2271:2264] ,data[2279:2272] ,data[2287:2280] ,data[2479:2472] ,data[2487:2480] ,data[2495:2488] ,data[2503:2496] ,data[2511:2504] ,data[2703:2696] ,data[2711:2704] ,data[2719:2712] ,data[2727:2720] ,data[2735:2728] };
end
284 :begin
 dPIn = {data[1815:1808] ,data[1823:1816] ,data[1831:1824] ,data[1839:1832] ,data[1847:1840] ,data[2039:2032] ,data[2047:2040] ,data[2055:2048] ,data[2063:2056] ,data[2071:2064] ,data[2263:2256] ,data[2271:2264] ,data[2279:2272] ,data[2287:2280] ,data[2295:2288] ,data[2487:2480] ,data[2495:2488] ,data[2503:2496] ,data[2511:2504] ,data[2519:2512] ,data[2711:2704] ,data[2719:2712] ,data[2727:2720] ,data[2735:2728] ,data[2743:2736] };
end
285 :begin
 dPIn = {data[1823:1816] ,data[1831:1824] ,data[1839:1832] ,data[1847:1840] ,data[1855:1848] ,data[2047:2040] ,data[2055:2048] ,data[2063:2056] ,data[2071:2064] ,data[2079:2072] ,data[2271:2264] ,data[2279:2272] ,data[2287:2280] ,data[2295:2288] ,data[2303:2296] ,data[2495:2488] ,data[2503:2496] ,data[2511:2504] ,data[2519:2512] ,data[2527:2520] ,data[2719:2712] ,data[2727:2720] ,data[2735:2728] ,data[2743:2736] ,data[2751:2744] };
end
286 :begin
 dPIn = {data[1831:1824] ,data[1839:1832] ,data[1847:1840] ,data[1855:1848] ,data[1863:1856] ,data[2055:2048] ,data[2063:2056] ,data[2071:2064] ,data[2079:2072] ,data[2087:2080] ,data[2279:2272] ,data[2287:2280] ,data[2295:2288] ,data[2303:2296] ,data[2311:2304] ,data[2503:2496] ,data[2511:2504] ,data[2519:2512] ,data[2527:2520] ,data[2535:2528] ,data[2727:2720] ,data[2735:2728] ,data[2743:2736] ,data[2751:2744] ,data[2759:2752] };
end
287 :begin
 dPIn = {data[1839:1832] ,data[1847:1840] ,data[1855:1848] ,data[1863:1856] ,data[1871:1864] ,data[2063:2056] ,data[2071:2064] ,data[2079:2072] ,data[2087:2080] ,data[2095:2088] ,data[2287:2280] ,data[2295:2288] ,data[2303:2296] ,data[2311:2304] ,data[2319:2312] ,data[2511:2504] ,data[2519:2512] ,data[2527:2520] ,data[2535:2528] ,data[2543:2536] ,data[2735:2728] ,data[2743:2736] ,data[2751:2744] ,data[2759:2752] ,data[2767:2760] };
end
288 :begin
 dPIn = {data[1847:1840] ,data[1855:1848] ,data[1863:1856] ,data[1871:1864] ,data[1879:1872] ,data[2071:2064] ,data[2079:2072] ,data[2087:2080] ,data[2095:2088] ,data[2103:2096] ,data[2295:2288] ,data[2303:2296] ,data[2311:2304] ,data[2319:2312] ,data[2327:2320] ,data[2519:2512] ,data[2527:2520] ,data[2535:2528] ,data[2543:2536] ,data[2551:2544] ,data[2743:2736] ,data[2751:2744] ,data[2759:2752] ,data[2767:2760] ,data[2775:2768] };
end
289 :begin
 dPIn = {data[1855:1848] ,data[1863:1856] ,data[1871:1864] ,data[1879:1872] ,data[1887:1880] ,data[2079:2072] ,data[2087:2080] ,data[2095:2088] ,data[2103:2096] ,data[2111:2104] ,data[2303:2296] ,data[2311:2304] ,data[2319:2312] ,data[2327:2320] ,data[2335:2328] ,data[2527:2520] ,data[2535:2528] ,data[2543:2536] ,data[2551:2544] ,data[2559:2552] ,data[2751:2744] ,data[2759:2752] ,data[2767:2760] ,data[2775:2768] ,data[2783:2776] };
end
290 :begin
 dPIn = {data[1863:1856] ,data[1871:1864] ,data[1879:1872] ,data[1887:1880] ,data[1895:1888] ,data[2087:2080] ,data[2095:2088] ,data[2103:2096] ,data[2111:2104] ,data[2119:2112] ,data[2311:2304] ,data[2319:2312] ,data[2327:2320] ,data[2335:2328] ,data[2343:2336] ,data[2535:2528] ,data[2543:2536] ,data[2551:2544] ,data[2559:2552] ,data[2567:2560] ,data[2759:2752] ,data[2767:2760] ,data[2775:2768] ,data[2783:2776] ,data[2791:2784] };
end
291 :begin
 dPIn = {data[1871:1864] ,data[1879:1872] ,data[1887:1880] ,data[1895:1888] ,data[1903:1896] ,data[2095:2088] ,data[2103:2096] ,data[2111:2104] ,data[2119:2112] ,data[2127:2120] ,data[2319:2312] ,data[2327:2320] ,data[2335:2328] ,data[2343:2336] ,data[2351:2344] ,data[2543:2536] ,data[2551:2544] ,data[2559:2552] ,data[2567:2560] ,data[2575:2568] ,data[2767:2760] ,data[2775:2768] ,data[2783:2776] ,data[2791:2784] ,data[2799:2792] };
end
292 :begin
 dPIn = {data[1879:1872] ,data[1887:1880] ,data[1895:1888] ,data[1903:1896] ,data[1911:1904] ,data[2103:2096] ,data[2111:2104] ,data[2119:2112] ,data[2127:2120] ,data[2135:2128] ,data[2327:2320] ,data[2335:2328] ,data[2343:2336] ,data[2351:2344] ,data[2359:2352] ,data[2551:2544] ,data[2559:2552] ,data[2567:2560] ,data[2575:2568] ,data[2583:2576] ,data[2775:2768] ,data[2783:2776] ,data[2791:2784] ,data[2799:2792] ,data[2807:2800] };
end
293 :begin
 dPIn = {data[1887:1880] ,data[1895:1888] ,data[1903:1896] ,data[1911:1904] ,data[1919:1912] ,data[2111:2104] ,data[2119:2112] ,data[2127:2120] ,data[2135:2128] ,data[2143:2136] ,data[2335:2328] ,data[2343:2336] ,data[2351:2344] ,data[2359:2352] ,data[2367:2360] ,data[2559:2552] ,data[2567:2560] ,data[2575:2568] ,data[2583:2576] ,data[2591:2584] ,data[2783:2776] ,data[2791:2784] ,data[2799:2792] ,data[2807:2800] ,data[2815:2808] };
end
294 :begin
 dPIn = {data[1895:1888] ,data[1903:1896] ,data[1911:1904] ,data[1919:1912] ,data[1927:1920] ,data[2119:2112] ,data[2127:2120] ,data[2135:2128] ,data[2143:2136] ,data[2151:2144] ,data[2343:2336] ,data[2351:2344] ,data[2359:2352] ,data[2367:2360] ,data[2375:2368] ,data[2567:2560] ,data[2575:2568] ,data[2583:2576] ,data[2591:2584] ,data[2599:2592] ,data[2791:2784] ,data[2799:2792] ,data[2807:2800] ,data[2815:2808] ,data[2823:2816] };
end
295 :begin
 dPIn = {data[1903:1896] ,data[1911:1904] ,data[1919:1912] ,data[1927:1920] ,data[1935:1928] ,data[2127:2120] ,data[2135:2128] ,data[2143:2136] ,data[2151:2144] ,data[2159:2152] ,data[2351:2344] ,data[2359:2352] ,data[2367:2360] ,data[2375:2368] ,data[2383:2376] ,data[2575:2568] ,data[2583:2576] ,data[2591:2584] ,data[2599:2592] ,data[2607:2600] ,data[2799:2792] ,data[2807:2800] ,data[2815:2808] ,data[2823:2816] ,data[2831:2824] };
end
296 :begin
 dPIn = {data[1911:1904] ,data[1919:1912] ,data[1927:1920] ,data[1935:1928] ,data[1943:1936] ,data[2135:2128] ,data[2143:2136] ,data[2151:2144] ,data[2159:2152] ,data[2167:2160] ,data[2359:2352] ,data[2367:2360] ,data[2375:2368] ,data[2383:2376] ,data[2391:2384] ,data[2583:2576] ,data[2591:2584] ,data[2599:2592] ,data[2607:2600] ,data[2615:2608] ,data[2807:2800] ,data[2815:2808] ,data[2823:2816] ,data[2831:2824] ,data[2839:2832] };
end
297 :begin
 dPIn = {data[1919:1912] ,data[1927:1920] ,data[1935:1928] ,data[1943:1936] ,data[1951:1944] ,data[2143:2136] ,data[2151:2144] ,data[2159:2152] ,data[2167:2160] ,data[2175:2168] ,data[2367:2360] ,data[2375:2368] ,data[2383:2376] ,data[2391:2384] ,data[2399:2392] ,data[2591:2584] ,data[2599:2592] ,data[2607:2600] ,data[2615:2608] ,data[2623:2616] ,data[2815:2808] ,data[2823:2816] ,data[2831:2824] ,data[2839:2832] ,data[2847:2840] };
end
298 :begin
 dPIn = {data[1927:1920] ,data[1935:1928] ,data[1943:1936] ,data[1951:1944] ,data[1959:1952] ,data[2151:2144] ,data[2159:2152] ,data[2167:2160] ,data[2175:2168] ,data[2183:2176] ,data[2375:2368] ,data[2383:2376] ,data[2391:2384] ,data[2399:2392] ,data[2407:2400] ,data[2599:2592] ,data[2607:2600] ,data[2615:2608] ,data[2623:2616] ,data[2631:2624] ,data[2823:2816] ,data[2831:2824] ,data[2839:2832] ,data[2847:2840] ,data[2855:2848] };
end
299 :begin
 dPIn = {data[1935:1928] ,data[1943:1936] ,data[1951:1944] ,data[1959:1952] ,data[1967:1960] ,data[2159:2152] ,data[2167:2160] ,data[2175:2168] ,data[2183:2176] ,data[2191:2184] ,data[2383:2376] ,data[2391:2384] ,data[2399:2392] ,data[2407:2400] ,data[2415:2408] ,data[2607:2600] ,data[2615:2608] ,data[2623:2616] ,data[2631:2624] ,data[2639:2632] ,data[2831:2824] ,data[2839:2832] ,data[2847:2840] ,data[2855:2848] ,data[2863:2856] };
end
300 :begin
 dPIn = {data[1943:1936] ,data[1951:1944] ,data[1959:1952] ,data[1967:1960] ,data[1975:1968] ,data[2167:2160] ,data[2175:2168] ,data[2183:2176] ,data[2191:2184] ,data[2199:2192] ,data[2391:2384] ,data[2399:2392] ,data[2407:2400] ,data[2415:2408] ,data[2423:2416] ,data[2615:2608] ,data[2623:2616] ,data[2631:2624] ,data[2639:2632] ,data[2647:2640] ,data[2839:2832] ,data[2847:2840] ,data[2855:2848] ,data[2863:2856] ,data[2871:2864] };
end
301 :begin
 dPIn = {data[1951:1944] ,data[1959:1952] ,data[1967:1960] ,data[1975:1968] ,data[1983:1976] ,data[2175:2168] ,data[2183:2176] ,data[2191:2184] ,data[2199:2192] ,data[2207:2200] ,data[2399:2392] ,data[2407:2400] ,data[2415:2408] ,data[2423:2416] ,data[2431:2424] ,data[2623:2616] ,data[2631:2624] ,data[2639:2632] ,data[2647:2640] ,data[2655:2648] ,data[2847:2840] ,data[2855:2848] ,data[2863:2856] ,data[2871:2864] ,data[2879:2872] };
end
302 :begin
 dPIn = {data[1959:1952] ,data[1967:1960] ,data[1975:1968] ,data[1983:1976] ,data[1991:1984] ,data[2183:2176] ,data[2191:2184] ,data[2199:2192] ,data[2207:2200] ,data[2215:2208] ,data[2407:2400] ,data[2415:2408] ,data[2423:2416] ,data[2431:2424] ,data[2439:2432] ,data[2631:2624] ,data[2639:2632] ,data[2647:2640] ,data[2655:2648] ,data[2663:2656] ,data[2855:2848] ,data[2863:2856] ,data[2871:2864] ,data[2879:2872] ,data[2887:2880] };
end
303 :begin
 dPIn = {data[1967:1960] ,data[1975:1968] ,data[1983:1976] ,data[1991:1984] ,data[1999:1992] ,data[2191:2184] ,data[2199:2192] ,data[2207:2200] ,data[2215:2208] ,data[2223:2216] ,data[2415:2408] ,data[2423:2416] ,data[2431:2424] ,data[2439:2432] ,data[2447:2440] ,data[2639:2632] ,data[2647:2640] ,data[2655:2648] ,data[2663:2656] ,data[2671:2664] ,data[2863:2856] ,data[2871:2864] ,data[2879:2872] ,data[2887:2880] ,data[2895:2888] };
end
304 :begin
 dPIn = {data[1975:1968] ,data[1983:1976] ,data[1991:1984] ,data[1999:1992] ,data[2007:2000] ,data[2199:2192] ,data[2207:2200] ,data[2215:2208] ,data[2223:2216] ,data[2231:2224] ,data[2423:2416] ,data[2431:2424] ,data[2439:2432] ,data[2447:2440] ,data[2455:2448] ,data[2647:2640] ,data[2655:2648] ,data[2663:2656] ,data[2671:2664] ,data[2679:2672] ,data[2871:2864] ,data[2879:2872] ,data[2887:2880] ,data[2895:2888] ,data[2903:2896] };
end
305 :begin
 dPIn = {data[1983:1976] ,data[1991:1984] ,data[1999:1992] ,data[2007:2000] ,data[2015:2008] ,data[2207:2200] ,data[2215:2208] ,data[2223:2216] ,data[2231:2224] ,data[2239:2232] ,data[2431:2424] ,data[2439:2432] ,data[2447:2440] ,data[2455:2448] ,data[2463:2456] ,data[2655:2648] ,data[2663:2656] ,data[2671:2664] ,data[2679:2672] ,data[2687:2680] ,data[2879:2872] ,data[2887:2880] ,data[2895:2888] ,data[2903:2896] ,data[2911:2904] };
end
306 :begin
 dPIn = {data[1991:1984] ,data[1999:1992] ,data[2007:2000] ,data[2015:2008] ,0 ,data[2215:2208] ,data[2223:2216] ,data[2231:2224] ,data[2239:2232] ,0 ,data[2439:2432] ,data[2447:2440] ,data[2455:2448] ,data[2463:2456] ,0 ,data[2663:2656] ,data[2671:2664] ,data[2679:2672] ,data[2687:2680] ,0 ,data[2887:2880] ,data[2895:2888] ,data[2903:2896] ,data[2911:2904] ,0 };
end
307 :begin
 dPIn = {data[1999:1992] ,data[2007:2000] ,data[2015:2008] ,0 ,0 ,data[2223:2216] ,data[2231:2224] ,data[2239:2232] ,0 ,0 ,data[2447:2440] ,data[2455:2448] ,data[2463:2456] ,0 ,0 ,data[2671:2664] ,data[2679:2672] ,data[2687:2680] ,0 ,0 ,data[2895:2888] ,data[2903:2896] ,data[2911:2904] ,0 ,0 };
end
308 :begin
 dPIn = {0 ,0 ,data[2023:2016] ,data[2031:2024] ,data[2039:2032] ,0 ,0 ,data[2247:2240] ,data[2255:2248] ,data[2263:2256] ,0 ,0 ,data[2471:2464] ,data[2479:2472] ,data[2487:2480] ,0 ,0 ,data[2695:2688] ,data[2703:2696] ,data[2711:2704] ,0 ,0 ,data[2919:2912] ,data[2927:2920] ,data[2935:2928] };
end
309 :begin
 dPIn = {0 ,data[2023:2016] ,data[2031:2024] ,data[2039:2032] ,data[2047:2040] ,0 ,data[2247:2240] ,data[2255:2248] ,data[2263:2256] ,data[2271:2264] ,0 ,data[2471:2464] ,data[2479:2472] ,data[2487:2480] ,data[2495:2488] ,0 ,data[2695:2688] ,data[2703:2696] ,data[2711:2704] ,data[2719:2712] ,0 ,data[2919:2912] ,data[2927:2920] ,data[2935:2928] ,data[2943:2936] };
end
310 :begin
 dPIn = {data[2023:2016] ,data[2031:2024] ,data[2039:2032] ,data[2047:2040] ,data[2055:2048] ,data[2247:2240] ,data[2255:2248] ,data[2263:2256] ,data[2271:2264] ,data[2279:2272] ,data[2471:2464] ,data[2479:2472] ,data[2487:2480] ,data[2495:2488] ,data[2503:2496] ,data[2695:2688] ,data[2703:2696] ,data[2711:2704] ,data[2719:2712] ,data[2727:2720] ,data[2919:2912] ,data[2927:2920] ,data[2935:2928] ,data[2943:2936] ,data[2951:2944] };
end
311 :begin
 dPIn = {data[2031:2024] ,data[2039:2032] ,data[2047:2040] ,data[2055:2048] ,data[2063:2056] ,data[2255:2248] ,data[2263:2256] ,data[2271:2264] ,data[2279:2272] ,data[2287:2280] ,data[2479:2472] ,data[2487:2480] ,data[2495:2488] ,data[2503:2496] ,data[2511:2504] ,data[2703:2696] ,data[2711:2704] ,data[2719:2712] ,data[2727:2720] ,data[2735:2728] ,data[2927:2920] ,data[2935:2928] ,data[2943:2936] ,data[2951:2944] ,data[2959:2952] };
end
312 :begin
 dPIn = {data[2039:2032] ,data[2047:2040] ,data[2055:2048] ,data[2063:2056] ,data[2071:2064] ,data[2263:2256] ,data[2271:2264] ,data[2279:2272] ,data[2287:2280] ,data[2295:2288] ,data[2487:2480] ,data[2495:2488] ,data[2503:2496] ,data[2511:2504] ,data[2519:2512] ,data[2711:2704] ,data[2719:2712] ,data[2727:2720] ,data[2735:2728] ,data[2743:2736] ,data[2935:2928] ,data[2943:2936] ,data[2951:2944] ,data[2959:2952] ,data[2967:2960] };
end
313 :begin
 dPIn = {data[2047:2040] ,data[2055:2048] ,data[2063:2056] ,data[2071:2064] ,data[2079:2072] ,data[2271:2264] ,data[2279:2272] ,data[2287:2280] ,data[2295:2288] ,data[2303:2296] ,data[2495:2488] ,data[2503:2496] ,data[2511:2504] ,data[2519:2512] ,data[2527:2520] ,data[2719:2712] ,data[2727:2720] ,data[2735:2728] ,data[2743:2736] ,data[2751:2744] ,data[2943:2936] ,data[2951:2944] ,data[2959:2952] ,data[2967:2960] ,data[2975:2968] };
end
314 :begin
 dPIn = {data[2055:2048] ,data[2063:2056] ,data[2071:2064] ,data[2079:2072] ,data[2087:2080] ,data[2279:2272] ,data[2287:2280] ,data[2295:2288] ,data[2303:2296] ,data[2311:2304] ,data[2503:2496] ,data[2511:2504] ,data[2519:2512] ,data[2527:2520] ,data[2535:2528] ,data[2727:2720] ,data[2735:2728] ,data[2743:2736] ,data[2751:2744] ,data[2759:2752] ,data[2951:2944] ,data[2959:2952] ,data[2967:2960] ,data[2975:2968] ,data[2983:2976] };
end
315 :begin
 dPIn = {data[2063:2056] ,data[2071:2064] ,data[2079:2072] ,data[2087:2080] ,data[2095:2088] ,data[2287:2280] ,data[2295:2288] ,data[2303:2296] ,data[2311:2304] ,data[2319:2312] ,data[2511:2504] ,data[2519:2512] ,data[2527:2520] ,data[2535:2528] ,data[2543:2536] ,data[2735:2728] ,data[2743:2736] ,data[2751:2744] ,data[2759:2752] ,data[2767:2760] ,data[2959:2952] ,data[2967:2960] ,data[2975:2968] ,data[2983:2976] ,data[2991:2984] };
end
316 :begin
 dPIn = {data[2071:2064] ,data[2079:2072] ,data[2087:2080] ,data[2095:2088] ,data[2103:2096] ,data[2295:2288] ,data[2303:2296] ,data[2311:2304] ,data[2319:2312] ,data[2327:2320] ,data[2519:2512] ,data[2527:2520] ,data[2535:2528] ,data[2543:2536] ,data[2551:2544] ,data[2743:2736] ,data[2751:2744] ,data[2759:2752] ,data[2767:2760] ,data[2775:2768] ,data[2967:2960] ,data[2975:2968] ,data[2983:2976] ,data[2991:2984] ,data[2999:2992] };
end
317 :begin
 dPIn = {data[2079:2072] ,data[2087:2080] ,data[2095:2088] ,data[2103:2096] ,data[2111:2104] ,data[2303:2296] ,data[2311:2304] ,data[2319:2312] ,data[2327:2320] ,data[2335:2328] ,data[2527:2520] ,data[2535:2528] ,data[2543:2536] ,data[2551:2544] ,data[2559:2552] ,data[2751:2744] ,data[2759:2752] ,data[2767:2760] ,data[2775:2768] ,data[2783:2776] ,data[2975:2968] ,data[2983:2976] ,data[2991:2984] ,data[2999:2992] ,data[3007:3000] };
end
318 :begin
 dPIn = {data[2087:2080] ,data[2095:2088] ,data[2103:2096] ,data[2111:2104] ,data[2119:2112] ,data[2311:2304] ,data[2319:2312] ,data[2327:2320] ,data[2335:2328] ,data[2343:2336] ,data[2535:2528] ,data[2543:2536] ,data[2551:2544] ,data[2559:2552] ,data[2567:2560] ,data[2759:2752] ,data[2767:2760] ,data[2775:2768] ,data[2783:2776] ,data[2791:2784] ,data[2983:2976] ,data[2991:2984] ,data[2999:2992] ,data[3007:3000] ,data[3015:3008] };
end
319 :begin
 dPIn = {data[2095:2088] ,data[2103:2096] ,data[2111:2104] ,data[2119:2112] ,data[2127:2120] ,data[2319:2312] ,data[2327:2320] ,data[2335:2328] ,data[2343:2336] ,data[2351:2344] ,data[2543:2536] ,data[2551:2544] ,data[2559:2552] ,data[2567:2560] ,data[2575:2568] ,data[2767:2760] ,data[2775:2768] ,data[2783:2776] ,data[2791:2784] ,data[2799:2792] ,data[2991:2984] ,data[2999:2992] ,data[3007:3000] ,data[3015:3008] ,data[3023:3016] };
end
320 :begin
 dPIn = {data[2103:2096] ,data[2111:2104] ,data[2119:2112] ,data[2127:2120] ,data[2135:2128] ,data[2327:2320] ,data[2335:2328] ,data[2343:2336] ,data[2351:2344] ,data[2359:2352] ,data[2551:2544] ,data[2559:2552] ,data[2567:2560] ,data[2575:2568] ,data[2583:2576] ,data[2775:2768] ,data[2783:2776] ,data[2791:2784] ,data[2799:2792] ,data[2807:2800] ,data[2999:2992] ,data[3007:3000] ,data[3015:3008] ,data[3023:3016] ,data[3031:3024] };
end
321 :begin
 dPIn = {data[2111:2104] ,data[2119:2112] ,data[2127:2120] ,data[2135:2128] ,data[2143:2136] ,data[2335:2328] ,data[2343:2336] ,data[2351:2344] ,data[2359:2352] ,data[2367:2360] ,data[2559:2552] ,data[2567:2560] ,data[2575:2568] ,data[2583:2576] ,data[2591:2584] ,data[2783:2776] ,data[2791:2784] ,data[2799:2792] ,data[2807:2800] ,data[2815:2808] ,data[3007:3000] ,data[3015:3008] ,data[3023:3016] ,data[3031:3024] ,data[3039:3032] };
end
322 :begin
 dPIn = {data[2119:2112] ,data[2127:2120] ,data[2135:2128] ,data[2143:2136] ,data[2151:2144] ,data[2343:2336] ,data[2351:2344] ,data[2359:2352] ,data[2367:2360] ,data[2375:2368] ,data[2567:2560] ,data[2575:2568] ,data[2583:2576] ,data[2591:2584] ,data[2599:2592] ,data[2791:2784] ,data[2799:2792] ,data[2807:2800] ,data[2815:2808] ,data[2823:2816] ,data[3015:3008] ,data[3023:3016] ,data[3031:3024] ,data[3039:3032] ,data[3047:3040] };
end
323 :begin
 dPIn = {data[2127:2120] ,data[2135:2128] ,data[2143:2136] ,data[2151:2144] ,data[2159:2152] ,data[2351:2344] ,data[2359:2352] ,data[2367:2360] ,data[2375:2368] ,data[2383:2376] ,data[2575:2568] ,data[2583:2576] ,data[2591:2584] ,data[2599:2592] ,data[2607:2600] ,data[2799:2792] ,data[2807:2800] ,data[2815:2808] ,data[2823:2816] ,data[2831:2824] ,data[3023:3016] ,data[3031:3024] ,data[3039:3032] ,data[3047:3040] ,data[3055:3048] };
end
324 :begin
 dPIn = {data[2135:2128] ,data[2143:2136] ,data[2151:2144] ,data[2159:2152] ,data[2167:2160] ,data[2359:2352] ,data[2367:2360] ,data[2375:2368] ,data[2383:2376] ,data[2391:2384] ,data[2583:2576] ,data[2591:2584] ,data[2599:2592] ,data[2607:2600] ,data[2615:2608] ,data[2807:2800] ,data[2815:2808] ,data[2823:2816] ,data[2831:2824] ,data[2839:2832] ,data[3031:3024] ,data[3039:3032] ,data[3047:3040] ,data[3055:3048] ,data[3063:3056] };
end
325 :begin
 dPIn = {data[2143:2136] ,data[2151:2144] ,data[2159:2152] ,data[2167:2160] ,data[2175:2168] ,data[2367:2360] ,data[2375:2368] ,data[2383:2376] ,data[2391:2384] ,data[2399:2392] ,data[2591:2584] ,data[2599:2592] ,data[2607:2600] ,data[2615:2608] ,data[2623:2616] ,data[2815:2808] ,data[2823:2816] ,data[2831:2824] ,data[2839:2832] ,data[2847:2840] ,data[3039:3032] ,data[3047:3040] ,data[3055:3048] ,data[3063:3056] ,data[3071:3064] };
end
326 :begin
 dPIn = {data[2151:2144] ,data[2159:2152] ,data[2167:2160] ,data[2175:2168] ,data[2183:2176] ,data[2375:2368] ,data[2383:2376] ,data[2391:2384] ,data[2399:2392] ,data[2407:2400] ,data[2599:2592] ,data[2607:2600] ,data[2615:2608] ,data[2623:2616] ,data[2631:2624] ,data[2823:2816] ,data[2831:2824] ,data[2839:2832] ,data[2847:2840] ,data[2855:2848] ,data[3047:3040] ,data[3055:3048] ,data[3063:3056] ,data[3071:3064] ,data[3079:3072] };
end
327 :begin
 dPIn = {data[2159:2152] ,data[2167:2160] ,data[2175:2168] ,data[2183:2176] ,data[2191:2184] ,data[2383:2376] ,data[2391:2384] ,data[2399:2392] ,data[2407:2400] ,data[2415:2408] ,data[2607:2600] ,data[2615:2608] ,data[2623:2616] ,data[2631:2624] ,data[2639:2632] ,data[2831:2824] ,data[2839:2832] ,data[2847:2840] ,data[2855:2848] ,data[2863:2856] ,data[3055:3048] ,data[3063:3056] ,data[3071:3064] ,data[3079:3072] ,data[3087:3080] };
end
328 :begin
 dPIn = {data[2167:2160] ,data[2175:2168] ,data[2183:2176] ,data[2191:2184] ,data[2199:2192] ,data[2391:2384] ,data[2399:2392] ,data[2407:2400] ,data[2415:2408] ,data[2423:2416] ,data[2615:2608] ,data[2623:2616] ,data[2631:2624] ,data[2639:2632] ,data[2647:2640] ,data[2839:2832] ,data[2847:2840] ,data[2855:2848] ,data[2863:2856] ,data[2871:2864] ,data[3063:3056] ,data[3071:3064] ,data[3079:3072] ,data[3087:3080] ,data[3095:3088] };
end
329 :begin
 dPIn = {data[2175:2168] ,data[2183:2176] ,data[2191:2184] ,data[2199:2192] ,data[2207:2200] ,data[2399:2392] ,data[2407:2400] ,data[2415:2408] ,data[2423:2416] ,data[2431:2424] ,data[2623:2616] ,data[2631:2624] ,data[2639:2632] ,data[2647:2640] ,data[2655:2648] ,data[2847:2840] ,data[2855:2848] ,data[2863:2856] ,data[2871:2864] ,data[2879:2872] ,data[3071:3064] ,data[3079:3072] ,data[3087:3080] ,data[3095:3088] ,data[3103:3096] };
end
330 :begin
 dPIn = {data[2183:2176] ,data[2191:2184] ,data[2199:2192] ,data[2207:2200] ,data[2215:2208] ,data[2407:2400] ,data[2415:2408] ,data[2423:2416] ,data[2431:2424] ,data[2439:2432] ,data[2631:2624] ,data[2639:2632] ,data[2647:2640] ,data[2655:2648] ,data[2663:2656] ,data[2855:2848] ,data[2863:2856] ,data[2871:2864] ,data[2879:2872] ,data[2887:2880] ,data[3079:3072] ,data[3087:3080] ,data[3095:3088] ,data[3103:3096] ,data[3111:3104] };
end
331 :begin
 dPIn = {data[2191:2184] ,data[2199:2192] ,data[2207:2200] ,data[2215:2208] ,data[2223:2216] ,data[2415:2408] ,data[2423:2416] ,data[2431:2424] ,data[2439:2432] ,data[2447:2440] ,data[2639:2632] ,data[2647:2640] ,data[2655:2648] ,data[2663:2656] ,data[2671:2664] ,data[2863:2856] ,data[2871:2864] ,data[2879:2872] ,data[2887:2880] ,data[2895:2888] ,data[3087:3080] ,data[3095:3088] ,data[3103:3096] ,data[3111:3104] ,data[3119:3112] };
end
332 :begin
 dPIn = {data[2199:2192] ,data[2207:2200] ,data[2215:2208] ,data[2223:2216] ,data[2231:2224] ,data[2423:2416] ,data[2431:2424] ,data[2439:2432] ,data[2447:2440] ,data[2455:2448] ,data[2647:2640] ,data[2655:2648] ,data[2663:2656] ,data[2671:2664] ,data[2679:2672] ,data[2871:2864] ,data[2879:2872] ,data[2887:2880] ,data[2895:2888] ,data[2903:2896] ,data[3095:3088] ,data[3103:3096] ,data[3111:3104] ,data[3119:3112] ,data[3127:3120] };
end
333 :begin
 dPIn = {data[2207:2200] ,data[2215:2208] ,data[2223:2216] ,data[2231:2224] ,data[2239:2232] ,data[2431:2424] ,data[2439:2432] ,data[2447:2440] ,data[2455:2448] ,data[2463:2456] ,data[2655:2648] ,data[2663:2656] ,data[2671:2664] ,data[2679:2672] ,data[2687:2680] ,data[2879:2872] ,data[2887:2880] ,data[2895:2888] ,data[2903:2896] ,data[2911:2904] ,data[3103:3096] ,data[3111:3104] ,data[3119:3112] ,data[3127:3120] ,data[3135:3128] };
end
334 :begin
 dPIn = {data[2215:2208] ,data[2223:2216] ,data[2231:2224] ,data[2239:2232] ,0 ,data[2439:2432] ,data[2447:2440] ,data[2455:2448] ,data[2463:2456] ,0 ,data[2663:2656] ,data[2671:2664] ,data[2679:2672] ,data[2687:2680] ,0 ,data[2887:2880] ,data[2895:2888] ,data[2903:2896] ,data[2911:2904] ,0 ,data[3111:3104] ,data[3119:3112] ,data[3127:3120] ,data[3135:3128] ,0 };
end
335 :begin
 dPIn = {data[2223:2216] ,data[2231:2224] ,data[2239:2232] ,0 ,0 ,data[2447:2440] ,data[2455:2448] ,data[2463:2456] ,0 ,0 ,data[2671:2664] ,data[2679:2672] ,data[2687:2680] ,0 ,0 ,data[2895:2888] ,data[2903:2896] ,data[2911:2904] ,0 ,0 ,data[3119:3112] ,data[3127:3120] ,data[3135:3128] ,0 ,0 };
end
336 :begin
 dPIn = {0 ,0 ,data[2247:2240] ,data[2255:2248] ,data[2263:2256] ,0 ,0 ,data[2471:2464] ,data[2479:2472] ,data[2487:2480] ,0 ,0 ,data[2695:2688] ,data[2703:2696] ,data[2711:2704] ,0 ,0 ,data[2919:2912] ,data[2927:2920] ,data[2935:2928] ,0 ,0 ,data[3143:3136] ,data[3151:3144] ,data[3159:3152] };
end
337 :begin
 dPIn = {0 ,data[2247:2240] ,data[2255:2248] ,data[2263:2256] ,data[2271:2264] ,0 ,data[2471:2464] ,data[2479:2472] ,data[2487:2480] ,data[2495:2488] ,0 ,data[2695:2688] ,data[2703:2696] ,data[2711:2704] ,data[2719:2712] ,0 ,data[2919:2912] ,data[2927:2920] ,data[2935:2928] ,data[2943:2936] ,0 ,data[3143:3136] ,data[3151:3144] ,data[3159:3152] ,data[3167:3160] };
end
338 :begin
 dPIn = {data[2247:2240] ,data[2255:2248] ,data[2263:2256] ,data[2271:2264] ,data[2279:2272] ,data[2471:2464] ,data[2479:2472] ,data[2487:2480] ,data[2495:2488] ,data[2503:2496] ,data[2695:2688] ,data[2703:2696] ,data[2711:2704] ,data[2719:2712] ,data[2727:2720] ,data[2919:2912] ,data[2927:2920] ,data[2935:2928] ,data[2943:2936] ,data[2951:2944] ,data[3143:3136] ,data[3151:3144] ,data[3159:3152] ,data[3167:3160] ,data[3175:3168] };
end
339 :begin
 dPIn = {data[2255:2248] ,data[2263:2256] ,data[2271:2264] ,data[2279:2272] ,data[2287:2280] ,data[2479:2472] ,data[2487:2480] ,data[2495:2488] ,data[2503:2496] ,data[2511:2504] ,data[2703:2696] ,data[2711:2704] ,data[2719:2712] ,data[2727:2720] ,data[2735:2728] ,data[2927:2920] ,data[2935:2928] ,data[2943:2936] ,data[2951:2944] ,data[2959:2952] ,data[3151:3144] ,data[3159:3152] ,data[3167:3160] ,data[3175:3168] ,data[3183:3176] };
end
340 :begin
 dPIn = {data[2263:2256] ,data[2271:2264] ,data[2279:2272] ,data[2287:2280] ,data[2295:2288] ,data[2487:2480] ,data[2495:2488] ,data[2503:2496] ,data[2511:2504] ,data[2519:2512] ,data[2711:2704] ,data[2719:2712] ,data[2727:2720] ,data[2735:2728] ,data[2743:2736] ,data[2935:2928] ,data[2943:2936] ,data[2951:2944] ,data[2959:2952] ,data[2967:2960] ,data[3159:3152] ,data[3167:3160] ,data[3175:3168] ,data[3183:3176] ,data[3191:3184] };
end
341 :begin
 dPIn = {data[2271:2264] ,data[2279:2272] ,data[2287:2280] ,data[2295:2288] ,data[2303:2296] ,data[2495:2488] ,data[2503:2496] ,data[2511:2504] ,data[2519:2512] ,data[2527:2520] ,data[2719:2712] ,data[2727:2720] ,data[2735:2728] ,data[2743:2736] ,data[2751:2744] ,data[2943:2936] ,data[2951:2944] ,data[2959:2952] ,data[2967:2960] ,data[2975:2968] ,data[3167:3160] ,data[3175:3168] ,data[3183:3176] ,data[3191:3184] ,data[3199:3192] };
end
342 :begin
 dPIn = {data[2279:2272] ,data[2287:2280] ,data[2295:2288] ,data[2303:2296] ,data[2311:2304] ,data[2503:2496] ,data[2511:2504] ,data[2519:2512] ,data[2527:2520] ,data[2535:2528] ,data[2727:2720] ,data[2735:2728] ,data[2743:2736] ,data[2751:2744] ,data[2759:2752] ,data[2951:2944] ,data[2959:2952] ,data[2967:2960] ,data[2975:2968] ,data[2983:2976] ,data[3175:3168] ,data[3183:3176] ,data[3191:3184] ,data[3199:3192] ,data[3207:3200] };
end
343 :begin
 dPIn = {data[2287:2280] ,data[2295:2288] ,data[2303:2296] ,data[2311:2304] ,data[2319:2312] ,data[2511:2504] ,data[2519:2512] ,data[2527:2520] ,data[2535:2528] ,data[2543:2536] ,data[2735:2728] ,data[2743:2736] ,data[2751:2744] ,data[2759:2752] ,data[2767:2760] ,data[2959:2952] ,data[2967:2960] ,data[2975:2968] ,data[2983:2976] ,data[2991:2984] ,data[3183:3176] ,data[3191:3184] ,data[3199:3192] ,data[3207:3200] ,data[3215:3208] };
end
344 :begin
 dPIn = {data[2295:2288] ,data[2303:2296] ,data[2311:2304] ,data[2319:2312] ,data[2327:2320] ,data[2519:2512] ,data[2527:2520] ,data[2535:2528] ,data[2543:2536] ,data[2551:2544] ,data[2743:2736] ,data[2751:2744] ,data[2759:2752] ,data[2767:2760] ,data[2775:2768] ,data[2967:2960] ,data[2975:2968] ,data[2983:2976] ,data[2991:2984] ,data[2999:2992] ,data[3191:3184] ,data[3199:3192] ,data[3207:3200] ,data[3215:3208] ,data[3223:3216] };
end
345 :begin
 dPIn = {data[2303:2296] ,data[2311:2304] ,data[2319:2312] ,data[2327:2320] ,data[2335:2328] ,data[2527:2520] ,data[2535:2528] ,data[2543:2536] ,data[2551:2544] ,data[2559:2552] ,data[2751:2744] ,data[2759:2752] ,data[2767:2760] ,data[2775:2768] ,data[2783:2776] ,data[2975:2968] ,data[2983:2976] ,data[2991:2984] ,data[2999:2992] ,data[3007:3000] ,data[3199:3192] ,data[3207:3200] ,data[3215:3208] ,data[3223:3216] ,data[3231:3224] };
end
346 :begin
 dPIn = {data[2311:2304] ,data[2319:2312] ,data[2327:2320] ,data[2335:2328] ,data[2343:2336] ,data[2535:2528] ,data[2543:2536] ,data[2551:2544] ,data[2559:2552] ,data[2567:2560] ,data[2759:2752] ,data[2767:2760] ,data[2775:2768] ,data[2783:2776] ,data[2791:2784] ,data[2983:2976] ,data[2991:2984] ,data[2999:2992] ,data[3007:3000] ,data[3015:3008] ,data[3207:3200] ,data[3215:3208] ,data[3223:3216] ,data[3231:3224] ,data[3239:3232] };
end
347 :begin
 dPIn = {data[2319:2312] ,data[2327:2320] ,data[2335:2328] ,data[2343:2336] ,data[2351:2344] ,data[2543:2536] ,data[2551:2544] ,data[2559:2552] ,data[2567:2560] ,data[2575:2568] ,data[2767:2760] ,data[2775:2768] ,data[2783:2776] ,data[2791:2784] ,data[2799:2792] ,data[2991:2984] ,data[2999:2992] ,data[3007:3000] ,data[3015:3008] ,data[3023:3016] ,data[3215:3208] ,data[3223:3216] ,data[3231:3224] ,data[3239:3232] ,data[3247:3240] };
end
348 :begin
 dPIn = {data[2327:2320] ,data[2335:2328] ,data[2343:2336] ,data[2351:2344] ,data[2359:2352] ,data[2551:2544] ,data[2559:2552] ,data[2567:2560] ,data[2575:2568] ,data[2583:2576] ,data[2775:2768] ,data[2783:2776] ,data[2791:2784] ,data[2799:2792] ,data[2807:2800] ,data[2999:2992] ,data[3007:3000] ,data[3015:3008] ,data[3023:3016] ,data[3031:3024] ,data[3223:3216] ,data[3231:3224] ,data[3239:3232] ,data[3247:3240] ,data[3255:3248] };
end
349 :begin
 dPIn = {data[2335:2328] ,data[2343:2336] ,data[2351:2344] ,data[2359:2352] ,data[2367:2360] ,data[2559:2552] ,data[2567:2560] ,data[2575:2568] ,data[2583:2576] ,data[2591:2584] ,data[2783:2776] ,data[2791:2784] ,data[2799:2792] ,data[2807:2800] ,data[2815:2808] ,data[3007:3000] ,data[3015:3008] ,data[3023:3016] ,data[3031:3024] ,data[3039:3032] ,data[3231:3224] ,data[3239:3232] ,data[3247:3240] ,data[3255:3248] ,data[3263:3256] };
end
350 :begin
 dPIn = {data[2343:2336] ,data[2351:2344] ,data[2359:2352] ,data[2367:2360] ,data[2375:2368] ,data[2567:2560] ,data[2575:2568] ,data[2583:2576] ,data[2591:2584] ,data[2599:2592] ,data[2791:2784] ,data[2799:2792] ,data[2807:2800] ,data[2815:2808] ,data[2823:2816] ,data[3015:3008] ,data[3023:3016] ,data[3031:3024] ,data[3039:3032] ,data[3047:3040] ,data[3239:3232] ,data[3247:3240] ,data[3255:3248] ,data[3263:3256] ,data[3271:3264] };
end
351 :begin
 dPIn = {data[2351:2344] ,data[2359:2352] ,data[2367:2360] ,data[2375:2368] ,data[2383:2376] ,data[2575:2568] ,data[2583:2576] ,data[2591:2584] ,data[2599:2592] ,data[2607:2600] ,data[2799:2792] ,data[2807:2800] ,data[2815:2808] ,data[2823:2816] ,data[2831:2824] ,data[3023:3016] ,data[3031:3024] ,data[3039:3032] ,data[3047:3040] ,data[3055:3048] ,data[3247:3240] ,data[3255:3248] ,data[3263:3256] ,data[3271:3264] ,data[3279:3272] };
end
352 :begin
 dPIn = {data[2359:2352] ,data[2367:2360] ,data[2375:2368] ,data[2383:2376] ,data[2391:2384] ,data[2583:2576] ,data[2591:2584] ,data[2599:2592] ,data[2607:2600] ,data[2615:2608] ,data[2807:2800] ,data[2815:2808] ,data[2823:2816] ,data[2831:2824] ,data[2839:2832] ,data[3031:3024] ,data[3039:3032] ,data[3047:3040] ,data[3055:3048] ,data[3063:3056] ,data[3255:3248] ,data[3263:3256] ,data[3271:3264] ,data[3279:3272] ,data[3287:3280] };
end
353 :begin
 dPIn = {data[2367:2360] ,data[2375:2368] ,data[2383:2376] ,data[2391:2384] ,data[2399:2392] ,data[2591:2584] ,data[2599:2592] ,data[2607:2600] ,data[2615:2608] ,data[2623:2616] ,data[2815:2808] ,data[2823:2816] ,data[2831:2824] ,data[2839:2832] ,data[2847:2840] ,data[3039:3032] ,data[3047:3040] ,data[3055:3048] ,data[3063:3056] ,data[3071:3064] ,data[3263:3256] ,data[3271:3264] ,data[3279:3272] ,data[3287:3280] ,data[3295:3288] };
end
354 :begin
 dPIn = {data[2375:2368] ,data[2383:2376] ,data[2391:2384] ,data[2399:2392] ,data[2407:2400] ,data[2599:2592] ,data[2607:2600] ,data[2615:2608] ,data[2623:2616] ,data[2631:2624] ,data[2823:2816] ,data[2831:2824] ,data[2839:2832] ,data[2847:2840] ,data[2855:2848] ,data[3047:3040] ,data[3055:3048] ,data[3063:3056] ,data[3071:3064] ,data[3079:3072] ,data[3271:3264] ,data[3279:3272] ,data[3287:3280] ,data[3295:3288] ,data[3303:3296] };
end
355 :begin
 dPIn = {data[2383:2376] ,data[2391:2384] ,data[2399:2392] ,data[2407:2400] ,data[2415:2408] ,data[2607:2600] ,data[2615:2608] ,data[2623:2616] ,data[2631:2624] ,data[2639:2632] ,data[2831:2824] ,data[2839:2832] ,data[2847:2840] ,data[2855:2848] ,data[2863:2856] ,data[3055:3048] ,data[3063:3056] ,data[3071:3064] ,data[3079:3072] ,data[3087:3080] ,data[3279:3272] ,data[3287:3280] ,data[3295:3288] ,data[3303:3296] ,data[3311:3304] };
end
356 :begin
 dPIn = {data[2391:2384] ,data[2399:2392] ,data[2407:2400] ,data[2415:2408] ,data[2423:2416] ,data[2615:2608] ,data[2623:2616] ,data[2631:2624] ,data[2639:2632] ,data[2647:2640] ,data[2839:2832] ,data[2847:2840] ,data[2855:2848] ,data[2863:2856] ,data[2871:2864] ,data[3063:3056] ,data[3071:3064] ,data[3079:3072] ,data[3087:3080] ,data[3095:3088] ,data[3287:3280] ,data[3295:3288] ,data[3303:3296] ,data[3311:3304] ,data[3319:3312] };
end
357 :begin
 dPIn = {data[2399:2392] ,data[2407:2400] ,data[2415:2408] ,data[2423:2416] ,data[2431:2424] ,data[2623:2616] ,data[2631:2624] ,data[2639:2632] ,data[2647:2640] ,data[2655:2648] ,data[2847:2840] ,data[2855:2848] ,data[2863:2856] ,data[2871:2864] ,data[2879:2872] ,data[3071:3064] ,data[3079:3072] ,data[3087:3080] ,data[3095:3088] ,data[3103:3096] ,data[3295:3288] ,data[3303:3296] ,data[3311:3304] ,data[3319:3312] ,data[3327:3320] };
end
358 :begin
 dPIn = {data[2407:2400] ,data[2415:2408] ,data[2423:2416] ,data[2431:2424] ,data[2439:2432] ,data[2631:2624] ,data[2639:2632] ,data[2647:2640] ,data[2655:2648] ,data[2663:2656] ,data[2855:2848] ,data[2863:2856] ,data[2871:2864] ,data[2879:2872] ,data[2887:2880] ,data[3079:3072] ,data[3087:3080] ,data[3095:3088] ,data[3103:3096] ,data[3111:3104] ,data[3303:3296] ,data[3311:3304] ,data[3319:3312] ,data[3327:3320] ,data[3335:3328] };
end
359 :begin
 dPIn = {data[2415:2408] ,data[2423:2416] ,data[2431:2424] ,data[2439:2432] ,data[2447:2440] ,data[2639:2632] ,data[2647:2640] ,data[2655:2648] ,data[2663:2656] ,data[2671:2664] ,data[2863:2856] ,data[2871:2864] ,data[2879:2872] ,data[2887:2880] ,data[2895:2888] ,data[3087:3080] ,data[3095:3088] ,data[3103:3096] ,data[3111:3104] ,data[3119:3112] ,data[3311:3304] ,data[3319:3312] ,data[3327:3320] ,data[3335:3328] ,data[3343:3336] };
end
360 :begin
 dPIn = {data[2423:2416] ,data[2431:2424] ,data[2439:2432] ,data[2447:2440] ,data[2455:2448] ,data[2647:2640] ,data[2655:2648] ,data[2663:2656] ,data[2671:2664] ,data[2679:2672] ,data[2871:2864] ,data[2879:2872] ,data[2887:2880] ,data[2895:2888] ,data[2903:2896] ,data[3095:3088] ,data[3103:3096] ,data[3111:3104] ,data[3119:3112] ,data[3127:3120] ,data[3319:3312] ,data[3327:3320] ,data[3335:3328] ,data[3343:3336] ,data[3351:3344] };
end
361 :begin
 dPIn = {data[2431:2424] ,data[2439:2432] ,data[2447:2440] ,data[2455:2448] ,data[2463:2456] ,data[2655:2648] ,data[2663:2656] ,data[2671:2664] ,data[2679:2672] ,data[2687:2680] ,data[2879:2872] ,data[2887:2880] ,data[2895:2888] ,data[2903:2896] ,data[2911:2904] ,data[3103:3096] ,data[3111:3104] ,data[3119:3112] ,data[3127:3120] ,data[3135:3128] ,data[3327:3320] ,data[3335:3328] ,data[3343:3336] ,data[3351:3344] ,data[3359:3352] };
end
362 :begin
 dPIn = {data[2439:2432] ,data[2447:2440] ,data[2455:2448] ,data[2463:2456] ,0 ,data[2663:2656] ,data[2671:2664] ,data[2679:2672] ,data[2687:2680] ,0 ,data[2887:2880] ,data[2895:2888] ,data[2903:2896] ,data[2911:2904] ,0 ,data[3111:3104] ,data[3119:3112] ,data[3127:3120] ,data[3135:3128] ,0 ,data[3335:3328] ,data[3343:3336] ,data[3351:3344] ,data[3359:3352] ,0 };
end
363 :begin
 dPIn = {data[2447:2440] ,data[2455:2448] ,data[2463:2456] ,0 ,0 ,data[2671:2664] ,data[2679:2672] ,data[2687:2680] ,0 ,0 ,data[2895:2888] ,data[2903:2896] ,data[2911:2904] ,0 ,0 ,data[3119:3112] ,data[3127:3120] ,data[3135:3128] ,0 ,0 ,data[3343:3336] ,data[3351:3344] ,data[3359:3352] ,0 ,0 };
end
364 :begin
 dPIn = {0 ,0 ,data[2471:2464] ,data[2479:2472] ,data[2487:2480] ,0 ,0 ,data[2695:2688] ,data[2703:2696] ,data[2711:2704] ,0 ,0 ,data[2919:2912] ,data[2927:2920] ,data[2935:2928] ,0 ,0 ,data[3143:3136] ,data[3151:3144] ,data[3159:3152] ,0 ,0 ,data[3367:3360] ,data[3375:3368] ,data[3383:3376] };
end
365 :begin
 dPIn = {0 ,data[2471:2464] ,data[2479:2472] ,data[2487:2480] ,data[2495:2488] ,0 ,data[2695:2688] ,data[2703:2696] ,data[2711:2704] ,data[2719:2712] ,0 ,data[2919:2912] ,data[2927:2920] ,data[2935:2928] ,data[2943:2936] ,0 ,data[3143:3136] ,data[3151:3144] ,data[3159:3152] ,data[3167:3160] ,0 ,data[3367:3360] ,data[3375:3368] ,data[3383:3376] ,data[3391:3384] };
end
366 :begin
 dPIn = {data[2471:2464] ,data[2479:2472] ,data[2487:2480] ,data[2495:2488] ,data[2503:2496] ,data[2695:2688] ,data[2703:2696] ,data[2711:2704] ,data[2719:2712] ,data[2727:2720] ,data[2919:2912] ,data[2927:2920] ,data[2935:2928] ,data[2943:2936] ,data[2951:2944] ,data[3143:3136] ,data[3151:3144] ,data[3159:3152] ,data[3167:3160] ,data[3175:3168] ,data[3367:3360] ,data[3375:3368] ,data[3383:3376] ,data[3391:3384] ,data[3399:3392] };
end
367 :begin
 dPIn = {data[2479:2472] ,data[2487:2480] ,data[2495:2488] ,data[2503:2496] ,data[2511:2504] ,data[2703:2696] ,data[2711:2704] ,data[2719:2712] ,data[2727:2720] ,data[2735:2728] ,data[2927:2920] ,data[2935:2928] ,data[2943:2936] ,data[2951:2944] ,data[2959:2952] ,data[3151:3144] ,data[3159:3152] ,data[3167:3160] ,data[3175:3168] ,data[3183:3176] ,data[3375:3368] ,data[3383:3376] ,data[3391:3384] ,data[3399:3392] ,data[3407:3400] };
end
368 :begin
 dPIn = {data[2487:2480] ,data[2495:2488] ,data[2503:2496] ,data[2511:2504] ,data[2519:2512] ,data[2711:2704] ,data[2719:2712] ,data[2727:2720] ,data[2735:2728] ,data[2743:2736] ,data[2935:2928] ,data[2943:2936] ,data[2951:2944] ,data[2959:2952] ,data[2967:2960] ,data[3159:3152] ,data[3167:3160] ,data[3175:3168] ,data[3183:3176] ,data[3191:3184] ,data[3383:3376] ,data[3391:3384] ,data[3399:3392] ,data[3407:3400] ,data[3415:3408] };
end
369 :begin
 dPIn = {data[2495:2488] ,data[2503:2496] ,data[2511:2504] ,data[2519:2512] ,data[2527:2520] ,data[2719:2712] ,data[2727:2720] ,data[2735:2728] ,data[2743:2736] ,data[2751:2744] ,data[2943:2936] ,data[2951:2944] ,data[2959:2952] ,data[2967:2960] ,data[2975:2968] ,data[3167:3160] ,data[3175:3168] ,data[3183:3176] ,data[3191:3184] ,data[3199:3192] ,data[3391:3384] ,data[3399:3392] ,data[3407:3400] ,data[3415:3408] ,data[3423:3416] };
end
370 :begin
 dPIn = {data[2503:2496] ,data[2511:2504] ,data[2519:2512] ,data[2527:2520] ,data[2535:2528] ,data[2727:2720] ,data[2735:2728] ,data[2743:2736] ,data[2751:2744] ,data[2759:2752] ,data[2951:2944] ,data[2959:2952] ,data[2967:2960] ,data[2975:2968] ,data[2983:2976] ,data[3175:3168] ,data[3183:3176] ,data[3191:3184] ,data[3199:3192] ,data[3207:3200] ,data[3399:3392] ,data[3407:3400] ,data[3415:3408] ,data[3423:3416] ,data[3431:3424] };
end
371 :begin
 dPIn = {data[2511:2504] ,data[2519:2512] ,data[2527:2520] ,data[2535:2528] ,data[2543:2536] ,data[2735:2728] ,data[2743:2736] ,data[2751:2744] ,data[2759:2752] ,data[2767:2760] ,data[2959:2952] ,data[2967:2960] ,data[2975:2968] ,data[2983:2976] ,data[2991:2984] ,data[3183:3176] ,data[3191:3184] ,data[3199:3192] ,data[3207:3200] ,data[3215:3208] ,data[3407:3400] ,data[3415:3408] ,data[3423:3416] ,data[3431:3424] ,data[3439:3432] };
end
372 :begin
 dPIn = {data[2519:2512] ,data[2527:2520] ,data[2535:2528] ,data[2543:2536] ,data[2551:2544] ,data[2743:2736] ,data[2751:2744] ,data[2759:2752] ,data[2767:2760] ,data[2775:2768] ,data[2967:2960] ,data[2975:2968] ,data[2983:2976] ,data[2991:2984] ,data[2999:2992] ,data[3191:3184] ,data[3199:3192] ,data[3207:3200] ,data[3215:3208] ,data[3223:3216] ,data[3415:3408] ,data[3423:3416] ,data[3431:3424] ,data[3439:3432] ,data[3447:3440] };
end
373 :begin
 dPIn = {data[2527:2520] ,data[2535:2528] ,data[2543:2536] ,data[2551:2544] ,data[2559:2552] ,data[2751:2744] ,data[2759:2752] ,data[2767:2760] ,data[2775:2768] ,data[2783:2776] ,data[2975:2968] ,data[2983:2976] ,data[2991:2984] ,data[2999:2992] ,data[3007:3000] ,data[3199:3192] ,data[3207:3200] ,data[3215:3208] ,data[3223:3216] ,data[3231:3224] ,data[3423:3416] ,data[3431:3424] ,data[3439:3432] ,data[3447:3440] ,data[3455:3448] };
end
374 :begin
 dPIn = {data[2535:2528] ,data[2543:2536] ,data[2551:2544] ,data[2559:2552] ,data[2567:2560] ,data[2759:2752] ,data[2767:2760] ,data[2775:2768] ,data[2783:2776] ,data[2791:2784] ,data[2983:2976] ,data[2991:2984] ,data[2999:2992] ,data[3007:3000] ,data[3015:3008] ,data[3207:3200] ,data[3215:3208] ,data[3223:3216] ,data[3231:3224] ,data[3239:3232] ,data[3431:3424] ,data[3439:3432] ,data[3447:3440] ,data[3455:3448] ,data[3463:3456] };
end
375 :begin
 dPIn = {data[2543:2536] ,data[2551:2544] ,data[2559:2552] ,data[2567:2560] ,data[2575:2568] ,data[2767:2760] ,data[2775:2768] ,data[2783:2776] ,data[2791:2784] ,data[2799:2792] ,data[2991:2984] ,data[2999:2992] ,data[3007:3000] ,data[3015:3008] ,data[3023:3016] ,data[3215:3208] ,data[3223:3216] ,data[3231:3224] ,data[3239:3232] ,data[3247:3240] ,data[3439:3432] ,data[3447:3440] ,data[3455:3448] ,data[3463:3456] ,data[3471:3464] };
end
376 :begin
 dPIn = {data[2551:2544] ,data[2559:2552] ,data[2567:2560] ,data[2575:2568] ,data[2583:2576] ,data[2775:2768] ,data[2783:2776] ,data[2791:2784] ,data[2799:2792] ,data[2807:2800] ,data[2999:2992] ,data[3007:3000] ,data[3015:3008] ,data[3023:3016] ,data[3031:3024] ,data[3223:3216] ,data[3231:3224] ,data[3239:3232] ,data[3247:3240] ,data[3255:3248] ,data[3447:3440] ,data[3455:3448] ,data[3463:3456] ,data[3471:3464] ,data[3479:3472] };
end
377 :begin
 dPIn = {data[2559:2552] ,data[2567:2560] ,data[2575:2568] ,data[2583:2576] ,data[2591:2584] ,data[2783:2776] ,data[2791:2784] ,data[2799:2792] ,data[2807:2800] ,data[2815:2808] ,data[3007:3000] ,data[3015:3008] ,data[3023:3016] ,data[3031:3024] ,data[3039:3032] ,data[3231:3224] ,data[3239:3232] ,data[3247:3240] ,data[3255:3248] ,data[3263:3256] ,data[3455:3448] ,data[3463:3456] ,data[3471:3464] ,data[3479:3472] ,data[3487:3480] };
end
378 :begin
 dPIn = {data[2567:2560] ,data[2575:2568] ,data[2583:2576] ,data[2591:2584] ,data[2599:2592] ,data[2791:2784] ,data[2799:2792] ,data[2807:2800] ,data[2815:2808] ,data[2823:2816] ,data[3015:3008] ,data[3023:3016] ,data[3031:3024] ,data[3039:3032] ,data[3047:3040] ,data[3239:3232] ,data[3247:3240] ,data[3255:3248] ,data[3263:3256] ,data[3271:3264] ,data[3463:3456] ,data[3471:3464] ,data[3479:3472] ,data[3487:3480] ,data[3495:3488] };
end
379 :begin
 dPIn = {data[2575:2568] ,data[2583:2576] ,data[2591:2584] ,data[2599:2592] ,data[2607:2600] ,data[2799:2792] ,data[2807:2800] ,data[2815:2808] ,data[2823:2816] ,data[2831:2824] ,data[3023:3016] ,data[3031:3024] ,data[3039:3032] ,data[3047:3040] ,data[3055:3048] ,data[3247:3240] ,data[3255:3248] ,data[3263:3256] ,data[3271:3264] ,data[3279:3272] ,data[3471:3464] ,data[3479:3472] ,data[3487:3480] ,data[3495:3488] ,data[3503:3496] };
end
380 :begin
 dPIn = {data[2583:2576] ,data[2591:2584] ,data[2599:2592] ,data[2607:2600] ,data[2615:2608] ,data[2807:2800] ,data[2815:2808] ,data[2823:2816] ,data[2831:2824] ,data[2839:2832] ,data[3031:3024] ,data[3039:3032] ,data[3047:3040] ,data[3055:3048] ,data[3063:3056] ,data[3255:3248] ,data[3263:3256] ,data[3271:3264] ,data[3279:3272] ,data[3287:3280] ,data[3479:3472] ,data[3487:3480] ,data[3495:3488] ,data[3503:3496] ,data[3511:3504] };
end
381 :begin
 dPIn = {data[2591:2584] ,data[2599:2592] ,data[2607:2600] ,data[2615:2608] ,data[2623:2616] ,data[2815:2808] ,data[2823:2816] ,data[2831:2824] ,data[2839:2832] ,data[2847:2840] ,data[3039:3032] ,data[3047:3040] ,data[3055:3048] ,data[3063:3056] ,data[3071:3064] ,data[3263:3256] ,data[3271:3264] ,data[3279:3272] ,data[3287:3280] ,data[3295:3288] ,data[3487:3480] ,data[3495:3488] ,data[3503:3496] ,data[3511:3504] ,data[3519:3512] };
end
382 :begin
 dPIn = {data[2599:2592] ,data[2607:2600] ,data[2615:2608] ,data[2623:2616] ,data[2631:2624] ,data[2823:2816] ,data[2831:2824] ,data[2839:2832] ,data[2847:2840] ,data[2855:2848] ,data[3047:3040] ,data[3055:3048] ,data[3063:3056] ,data[3071:3064] ,data[3079:3072] ,data[3271:3264] ,data[3279:3272] ,data[3287:3280] ,data[3295:3288] ,data[3303:3296] ,data[3495:3488] ,data[3503:3496] ,data[3511:3504] ,data[3519:3512] ,data[3527:3520] };
end
383 :begin
 dPIn = {data[2607:2600] ,data[2615:2608] ,data[2623:2616] ,data[2631:2624] ,data[2639:2632] ,data[2831:2824] ,data[2839:2832] ,data[2847:2840] ,data[2855:2848] ,data[2863:2856] ,data[3055:3048] ,data[3063:3056] ,data[3071:3064] ,data[3079:3072] ,data[3087:3080] ,data[3279:3272] ,data[3287:3280] ,data[3295:3288] ,data[3303:3296] ,data[3311:3304] ,data[3503:3496] ,data[3511:3504] ,data[3519:3512] ,data[3527:3520] ,data[3535:3528] };
end
384 :begin
 dPIn = {data[2615:2608] ,data[2623:2616] ,data[2631:2624] ,data[2639:2632] ,data[2647:2640] ,data[2839:2832] ,data[2847:2840] ,data[2855:2848] ,data[2863:2856] ,data[2871:2864] ,data[3063:3056] ,data[3071:3064] ,data[3079:3072] ,data[3087:3080] ,data[3095:3088] ,data[3287:3280] ,data[3295:3288] ,data[3303:3296] ,data[3311:3304] ,data[3319:3312] ,data[3511:3504] ,data[3519:3512] ,data[3527:3520] ,data[3535:3528] ,data[3543:3536] };
end
385 :begin
 dPIn = {data[2623:2616] ,data[2631:2624] ,data[2639:2632] ,data[2647:2640] ,data[2655:2648] ,data[2847:2840] ,data[2855:2848] ,data[2863:2856] ,data[2871:2864] ,data[2879:2872] ,data[3071:3064] ,data[3079:3072] ,data[3087:3080] ,data[3095:3088] ,data[3103:3096] ,data[3295:3288] ,data[3303:3296] ,data[3311:3304] ,data[3319:3312] ,data[3327:3320] ,data[3519:3512] ,data[3527:3520] ,data[3535:3528] ,data[3543:3536] ,data[3551:3544] };
end
386 :begin
 dPIn = {data[2631:2624] ,data[2639:2632] ,data[2647:2640] ,data[2655:2648] ,data[2663:2656] ,data[2855:2848] ,data[2863:2856] ,data[2871:2864] ,data[2879:2872] ,data[2887:2880] ,data[3079:3072] ,data[3087:3080] ,data[3095:3088] ,data[3103:3096] ,data[3111:3104] ,data[3303:3296] ,data[3311:3304] ,data[3319:3312] ,data[3327:3320] ,data[3335:3328] ,data[3527:3520] ,data[3535:3528] ,data[3543:3536] ,data[3551:3544] ,data[3559:3552] };
end
387 :begin
 dPIn = {data[2639:2632] ,data[2647:2640] ,data[2655:2648] ,data[2663:2656] ,data[2671:2664] ,data[2863:2856] ,data[2871:2864] ,data[2879:2872] ,data[2887:2880] ,data[2895:2888] ,data[3087:3080] ,data[3095:3088] ,data[3103:3096] ,data[3111:3104] ,data[3119:3112] ,data[3311:3304] ,data[3319:3312] ,data[3327:3320] ,data[3335:3328] ,data[3343:3336] ,data[3535:3528] ,data[3543:3536] ,data[3551:3544] ,data[3559:3552] ,data[3567:3560] };
end
388 :begin
 dPIn = {data[2647:2640] ,data[2655:2648] ,data[2663:2656] ,data[2671:2664] ,data[2679:2672] ,data[2871:2864] ,data[2879:2872] ,data[2887:2880] ,data[2895:2888] ,data[2903:2896] ,data[3095:3088] ,data[3103:3096] ,data[3111:3104] ,data[3119:3112] ,data[3127:3120] ,data[3319:3312] ,data[3327:3320] ,data[3335:3328] ,data[3343:3336] ,data[3351:3344] ,data[3543:3536] ,data[3551:3544] ,data[3559:3552] ,data[3567:3560] ,data[3575:3568] };
end
389 :begin
 dPIn = {data[2655:2648] ,data[2663:2656] ,data[2671:2664] ,data[2679:2672] ,data[2687:2680] ,data[2879:2872] ,data[2887:2880] ,data[2895:2888] ,data[2903:2896] ,data[2911:2904] ,data[3103:3096] ,data[3111:3104] ,data[3119:3112] ,data[3127:3120] ,data[3135:3128] ,data[3327:3320] ,data[3335:3328] ,data[3343:3336] ,data[3351:3344] ,data[3359:3352] ,data[3551:3544] ,data[3559:3552] ,data[3567:3560] ,data[3575:3568] ,data[3583:3576] };
end
390 :begin
 dPIn = {data[2663:2656] ,data[2671:2664] ,data[2679:2672] ,data[2687:2680] ,0 ,data[2887:2880] ,data[2895:2888] ,data[2903:2896] ,data[2911:2904] ,0 ,data[3111:3104] ,data[3119:3112] ,data[3127:3120] ,data[3135:3128] ,0 ,data[3335:3328] ,data[3343:3336] ,data[3351:3344] ,data[3359:3352] ,0 ,data[3559:3552] ,data[3567:3560] ,data[3575:3568] ,data[3583:3576] ,0 };
end
391 :begin
 dPIn = {data[2671:2664] ,data[2679:2672] ,data[2687:2680] ,0 ,0 ,data[2895:2888] ,data[2903:2896] ,data[2911:2904] ,0 ,0 ,data[3119:3112] ,data[3127:3120] ,data[3135:3128] ,0 ,0 ,data[3343:3336] ,data[3351:3344] ,data[3359:3352] ,0 ,0 ,data[3567:3560] ,data[3575:3568] ,data[3583:3576] ,0 ,0 };
end
392 :begin
 dPIn = {0 ,0 ,data[2695:2688] ,data[2703:2696] ,data[2711:2704] ,0 ,0 ,data[2919:2912] ,data[2927:2920] ,data[2935:2928] ,0 ,0 ,data[3143:3136] ,data[3151:3144] ,data[3159:3152] ,0 ,0 ,data[3367:3360] ,data[3375:3368] ,data[3383:3376] ,0 ,0 ,data[3591:3584] ,data[3599:3592] ,data[3607:3600] };
end
393 :begin
 dPIn = {0 ,data[2695:2688] ,data[2703:2696] ,data[2711:2704] ,data[2719:2712] ,0 ,data[2919:2912] ,data[2927:2920] ,data[2935:2928] ,data[2943:2936] ,0 ,data[3143:3136] ,data[3151:3144] ,data[3159:3152] ,data[3167:3160] ,0 ,data[3367:3360] ,data[3375:3368] ,data[3383:3376] ,data[3391:3384] ,0 ,data[3591:3584] ,data[3599:3592] ,data[3607:3600] ,data[3615:3608] };
end
394 :begin
 dPIn = {data[2695:2688] ,data[2703:2696] ,data[2711:2704] ,data[2719:2712] ,data[2727:2720] ,data[2919:2912] ,data[2927:2920] ,data[2935:2928] ,data[2943:2936] ,data[2951:2944] ,data[3143:3136] ,data[3151:3144] ,data[3159:3152] ,data[3167:3160] ,data[3175:3168] ,data[3367:3360] ,data[3375:3368] ,data[3383:3376] ,data[3391:3384] ,data[3399:3392] ,data[3591:3584] ,data[3599:3592] ,data[3607:3600] ,data[3615:3608] ,data[3623:3616] };
end
395 :begin
 dPIn = {data[2703:2696] ,data[2711:2704] ,data[2719:2712] ,data[2727:2720] ,data[2735:2728] ,data[2927:2920] ,data[2935:2928] ,data[2943:2936] ,data[2951:2944] ,data[2959:2952] ,data[3151:3144] ,data[3159:3152] ,data[3167:3160] ,data[3175:3168] ,data[3183:3176] ,data[3375:3368] ,data[3383:3376] ,data[3391:3384] ,data[3399:3392] ,data[3407:3400] ,data[3599:3592] ,data[3607:3600] ,data[3615:3608] ,data[3623:3616] ,data[3631:3624] };
end
396 :begin
 dPIn = {data[2711:2704] ,data[2719:2712] ,data[2727:2720] ,data[2735:2728] ,data[2743:2736] ,data[2935:2928] ,data[2943:2936] ,data[2951:2944] ,data[2959:2952] ,data[2967:2960] ,data[3159:3152] ,data[3167:3160] ,data[3175:3168] ,data[3183:3176] ,data[3191:3184] ,data[3383:3376] ,data[3391:3384] ,data[3399:3392] ,data[3407:3400] ,data[3415:3408] ,data[3607:3600] ,data[3615:3608] ,data[3623:3616] ,data[3631:3624] ,data[3639:3632] };
end
397 :begin
 dPIn = {data[2719:2712] ,data[2727:2720] ,data[2735:2728] ,data[2743:2736] ,data[2751:2744] ,data[2943:2936] ,data[2951:2944] ,data[2959:2952] ,data[2967:2960] ,data[2975:2968] ,data[3167:3160] ,data[3175:3168] ,data[3183:3176] ,data[3191:3184] ,data[3199:3192] ,data[3391:3384] ,data[3399:3392] ,data[3407:3400] ,data[3415:3408] ,data[3423:3416] ,data[3615:3608] ,data[3623:3616] ,data[3631:3624] ,data[3639:3632] ,data[3647:3640] };
end
398 :begin
 dPIn = {data[2727:2720] ,data[2735:2728] ,data[2743:2736] ,data[2751:2744] ,data[2759:2752] ,data[2951:2944] ,data[2959:2952] ,data[2967:2960] ,data[2975:2968] ,data[2983:2976] ,data[3175:3168] ,data[3183:3176] ,data[3191:3184] ,data[3199:3192] ,data[3207:3200] ,data[3399:3392] ,data[3407:3400] ,data[3415:3408] ,data[3423:3416] ,data[3431:3424] ,data[3623:3616] ,data[3631:3624] ,data[3639:3632] ,data[3647:3640] ,data[3655:3648] };
end
399 :begin
 dPIn = {data[2735:2728] ,data[2743:2736] ,data[2751:2744] ,data[2759:2752] ,data[2767:2760] ,data[2959:2952] ,data[2967:2960] ,data[2975:2968] ,data[2983:2976] ,data[2991:2984] ,data[3183:3176] ,data[3191:3184] ,data[3199:3192] ,data[3207:3200] ,data[3215:3208] ,data[3407:3400] ,data[3415:3408] ,data[3423:3416] ,data[3431:3424] ,data[3439:3432] ,data[3631:3624] ,data[3639:3632] ,data[3647:3640] ,data[3655:3648] ,data[3663:3656] };
end
400 :begin
 dPIn = {data[2743:2736] ,data[2751:2744] ,data[2759:2752] ,data[2767:2760] ,data[2775:2768] ,data[2967:2960] ,data[2975:2968] ,data[2983:2976] ,data[2991:2984] ,data[2999:2992] ,data[3191:3184] ,data[3199:3192] ,data[3207:3200] ,data[3215:3208] ,data[3223:3216] ,data[3415:3408] ,data[3423:3416] ,data[3431:3424] ,data[3439:3432] ,data[3447:3440] ,data[3639:3632] ,data[3647:3640] ,data[3655:3648] ,data[3663:3656] ,data[3671:3664] };
end
401 :begin
 dPIn = {data[2751:2744] ,data[2759:2752] ,data[2767:2760] ,data[2775:2768] ,data[2783:2776] ,data[2975:2968] ,data[2983:2976] ,data[2991:2984] ,data[2999:2992] ,data[3007:3000] ,data[3199:3192] ,data[3207:3200] ,data[3215:3208] ,data[3223:3216] ,data[3231:3224] ,data[3423:3416] ,data[3431:3424] ,data[3439:3432] ,data[3447:3440] ,data[3455:3448] ,data[3647:3640] ,data[3655:3648] ,data[3663:3656] ,data[3671:3664] ,data[3679:3672] };
end
402 :begin
 dPIn = {data[2759:2752] ,data[2767:2760] ,data[2775:2768] ,data[2783:2776] ,data[2791:2784] ,data[2983:2976] ,data[2991:2984] ,data[2999:2992] ,data[3007:3000] ,data[3015:3008] ,data[3207:3200] ,data[3215:3208] ,data[3223:3216] ,data[3231:3224] ,data[3239:3232] ,data[3431:3424] ,data[3439:3432] ,data[3447:3440] ,data[3455:3448] ,data[3463:3456] ,data[3655:3648] ,data[3663:3656] ,data[3671:3664] ,data[3679:3672] ,data[3687:3680] };
end
403 :begin
 dPIn = {data[2767:2760] ,data[2775:2768] ,data[2783:2776] ,data[2791:2784] ,data[2799:2792] ,data[2991:2984] ,data[2999:2992] ,data[3007:3000] ,data[3015:3008] ,data[3023:3016] ,data[3215:3208] ,data[3223:3216] ,data[3231:3224] ,data[3239:3232] ,data[3247:3240] ,data[3439:3432] ,data[3447:3440] ,data[3455:3448] ,data[3463:3456] ,data[3471:3464] ,data[3663:3656] ,data[3671:3664] ,data[3679:3672] ,data[3687:3680] ,data[3695:3688] };
end
404 :begin
 dPIn = {data[2775:2768] ,data[2783:2776] ,data[2791:2784] ,data[2799:2792] ,data[2807:2800] ,data[2999:2992] ,data[3007:3000] ,data[3015:3008] ,data[3023:3016] ,data[3031:3024] ,data[3223:3216] ,data[3231:3224] ,data[3239:3232] ,data[3247:3240] ,data[3255:3248] ,data[3447:3440] ,data[3455:3448] ,data[3463:3456] ,data[3471:3464] ,data[3479:3472] ,data[3671:3664] ,data[3679:3672] ,data[3687:3680] ,data[3695:3688] ,data[3703:3696] };
end
405 :begin
 dPIn = {data[2783:2776] ,data[2791:2784] ,data[2799:2792] ,data[2807:2800] ,data[2815:2808] ,data[3007:3000] ,data[3015:3008] ,data[3023:3016] ,data[3031:3024] ,data[3039:3032] ,data[3231:3224] ,data[3239:3232] ,data[3247:3240] ,data[3255:3248] ,data[3263:3256] ,data[3455:3448] ,data[3463:3456] ,data[3471:3464] ,data[3479:3472] ,data[3487:3480] ,data[3679:3672] ,data[3687:3680] ,data[3695:3688] ,data[3703:3696] ,data[3711:3704] };
end
406 :begin
 dPIn = {data[2791:2784] ,data[2799:2792] ,data[2807:2800] ,data[2815:2808] ,data[2823:2816] ,data[3015:3008] ,data[3023:3016] ,data[3031:3024] ,data[3039:3032] ,data[3047:3040] ,data[3239:3232] ,data[3247:3240] ,data[3255:3248] ,data[3263:3256] ,data[3271:3264] ,data[3463:3456] ,data[3471:3464] ,data[3479:3472] ,data[3487:3480] ,data[3495:3488] ,data[3687:3680] ,data[3695:3688] ,data[3703:3696] ,data[3711:3704] ,data[3719:3712] };
end
407 :begin
 dPIn = {data[2799:2792] ,data[2807:2800] ,data[2815:2808] ,data[2823:2816] ,data[2831:2824] ,data[3023:3016] ,data[3031:3024] ,data[3039:3032] ,data[3047:3040] ,data[3055:3048] ,data[3247:3240] ,data[3255:3248] ,data[3263:3256] ,data[3271:3264] ,data[3279:3272] ,data[3471:3464] ,data[3479:3472] ,data[3487:3480] ,data[3495:3488] ,data[3503:3496] ,data[3695:3688] ,data[3703:3696] ,data[3711:3704] ,data[3719:3712] ,data[3727:3720] };
end
408 :begin
 dPIn = {data[2807:2800] ,data[2815:2808] ,data[2823:2816] ,data[2831:2824] ,data[2839:2832] ,data[3031:3024] ,data[3039:3032] ,data[3047:3040] ,data[3055:3048] ,data[3063:3056] ,data[3255:3248] ,data[3263:3256] ,data[3271:3264] ,data[3279:3272] ,data[3287:3280] ,data[3479:3472] ,data[3487:3480] ,data[3495:3488] ,data[3503:3496] ,data[3511:3504] ,data[3703:3696] ,data[3711:3704] ,data[3719:3712] ,data[3727:3720] ,data[3735:3728] };
end
409 :begin
 dPIn = {data[2815:2808] ,data[2823:2816] ,data[2831:2824] ,data[2839:2832] ,data[2847:2840] ,data[3039:3032] ,data[3047:3040] ,data[3055:3048] ,data[3063:3056] ,data[3071:3064] ,data[3263:3256] ,data[3271:3264] ,data[3279:3272] ,data[3287:3280] ,data[3295:3288] ,data[3487:3480] ,data[3495:3488] ,data[3503:3496] ,data[3511:3504] ,data[3519:3512] ,data[3711:3704] ,data[3719:3712] ,data[3727:3720] ,data[3735:3728] ,data[3743:3736] };
end
410 :begin
 dPIn = {data[2823:2816] ,data[2831:2824] ,data[2839:2832] ,data[2847:2840] ,data[2855:2848] ,data[3047:3040] ,data[3055:3048] ,data[3063:3056] ,data[3071:3064] ,data[3079:3072] ,data[3271:3264] ,data[3279:3272] ,data[3287:3280] ,data[3295:3288] ,data[3303:3296] ,data[3495:3488] ,data[3503:3496] ,data[3511:3504] ,data[3519:3512] ,data[3527:3520] ,data[3719:3712] ,data[3727:3720] ,data[3735:3728] ,data[3743:3736] ,data[3751:3744] };
end
411 :begin
 dPIn = {data[2831:2824] ,data[2839:2832] ,data[2847:2840] ,data[2855:2848] ,data[2863:2856] ,data[3055:3048] ,data[3063:3056] ,data[3071:3064] ,data[3079:3072] ,data[3087:3080] ,data[3279:3272] ,data[3287:3280] ,data[3295:3288] ,data[3303:3296] ,data[3311:3304] ,data[3503:3496] ,data[3511:3504] ,data[3519:3512] ,data[3527:3520] ,data[3535:3528] ,data[3727:3720] ,data[3735:3728] ,data[3743:3736] ,data[3751:3744] ,data[3759:3752] };
end
412 :begin
 dPIn = {data[2839:2832] ,data[2847:2840] ,data[2855:2848] ,data[2863:2856] ,data[2871:2864] ,data[3063:3056] ,data[3071:3064] ,data[3079:3072] ,data[3087:3080] ,data[3095:3088] ,data[3287:3280] ,data[3295:3288] ,data[3303:3296] ,data[3311:3304] ,data[3319:3312] ,data[3511:3504] ,data[3519:3512] ,data[3527:3520] ,data[3535:3528] ,data[3543:3536] ,data[3735:3728] ,data[3743:3736] ,data[3751:3744] ,data[3759:3752] ,data[3767:3760] };
end
413 :begin
 dPIn = {data[2847:2840] ,data[2855:2848] ,data[2863:2856] ,data[2871:2864] ,data[2879:2872] ,data[3071:3064] ,data[3079:3072] ,data[3087:3080] ,data[3095:3088] ,data[3103:3096] ,data[3295:3288] ,data[3303:3296] ,data[3311:3304] ,data[3319:3312] ,data[3327:3320] ,data[3519:3512] ,data[3527:3520] ,data[3535:3528] ,data[3543:3536] ,data[3551:3544] ,data[3743:3736] ,data[3751:3744] ,data[3759:3752] ,data[3767:3760] ,data[3775:3768] };
end
414 :begin
 dPIn = {data[2855:2848] ,data[2863:2856] ,data[2871:2864] ,data[2879:2872] ,data[2887:2880] ,data[3079:3072] ,data[3087:3080] ,data[3095:3088] ,data[3103:3096] ,data[3111:3104] ,data[3303:3296] ,data[3311:3304] ,data[3319:3312] ,data[3327:3320] ,data[3335:3328] ,data[3527:3520] ,data[3535:3528] ,data[3543:3536] ,data[3551:3544] ,data[3559:3552] ,data[3751:3744] ,data[3759:3752] ,data[3767:3760] ,data[3775:3768] ,data[3783:3776] };
end
415 :begin
 dPIn = {data[2863:2856] ,data[2871:2864] ,data[2879:2872] ,data[2887:2880] ,data[2895:2888] ,data[3087:3080] ,data[3095:3088] ,data[3103:3096] ,data[3111:3104] ,data[3119:3112] ,data[3311:3304] ,data[3319:3312] ,data[3327:3320] ,data[3335:3328] ,data[3343:3336] ,data[3535:3528] ,data[3543:3536] ,data[3551:3544] ,data[3559:3552] ,data[3567:3560] ,data[3759:3752] ,data[3767:3760] ,data[3775:3768] ,data[3783:3776] ,data[3791:3784] };
end
416 :begin
 dPIn = {data[2871:2864] ,data[2879:2872] ,data[2887:2880] ,data[2895:2888] ,data[2903:2896] ,data[3095:3088] ,data[3103:3096] ,data[3111:3104] ,data[3119:3112] ,data[3127:3120] ,data[3319:3312] ,data[3327:3320] ,data[3335:3328] ,data[3343:3336] ,data[3351:3344] ,data[3543:3536] ,data[3551:3544] ,data[3559:3552] ,data[3567:3560] ,data[3575:3568] ,data[3767:3760] ,data[3775:3768] ,data[3783:3776] ,data[3791:3784] ,data[3799:3792] };
end
417 :begin
 dPIn = {data[2879:2872] ,data[2887:2880] ,data[2895:2888] ,data[2903:2896] ,data[2911:2904] ,data[3103:3096] ,data[3111:3104] ,data[3119:3112] ,data[3127:3120] ,data[3135:3128] ,data[3327:3320] ,data[3335:3328] ,data[3343:3336] ,data[3351:3344] ,data[3359:3352] ,data[3551:3544] ,data[3559:3552] ,data[3567:3560] ,data[3575:3568] ,data[3583:3576] ,data[3775:3768] ,data[3783:3776] ,data[3791:3784] ,data[3799:3792] ,data[3807:3800] };
end
418 :begin
 dPIn = {data[2887:2880] ,data[2895:2888] ,data[2903:2896] ,data[2911:2904] ,0 ,data[3111:3104] ,data[3119:3112] ,data[3127:3120] ,data[3135:3128] ,0 ,data[3335:3328] ,data[3343:3336] ,data[3351:3344] ,data[3359:3352] ,0 ,data[3559:3552] ,data[3567:3560] ,data[3575:3568] ,data[3583:3576] ,0 ,data[3783:3776] ,data[3791:3784] ,data[3799:3792] ,data[3807:3800] ,0 };
end
419 :begin
 dPIn = {data[2895:2888] ,data[2903:2896] ,data[2911:2904] ,0 ,0 ,data[3119:3112] ,data[3127:3120] ,data[3135:3128] ,0 ,0 ,data[3343:3336] ,data[3351:3344] ,data[3359:3352] ,0 ,0 ,data[3567:3560] ,data[3575:3568] ,data[3583:3576] ,0 ,0 ,data[3791:3784] ,data[3799:3792] ,data[3807:3800] ,0 ,0 };
end
420 :begin
 dPIn = {0 ,0 ,data[2919:2912] ,data[2927:2920] ,data[2935:2928] ,0 ,0 ,data[3143:3136] ,data[3151:3144] ,data[3159:3152] ,0 ,0 ,data[3367:3360] ,data[3375:3368] ,data[3383:3376] ,0 ,0 ,data[3591:3584] ,data[3599:3592] ,data[3607:3600] ,0 ,0 ,data[3815:3808] ,data[3823:3816] ,data[3831:3824] };
end
421 :begin
 dPIn = {0 ,data[2919:2912] ,data[2927:2920] ,data[2935:2928] ,data[2943:2936] ,0 ,data[3143:3136] ,data[3151:3144] ,data[3159:3152] ,data[3167:3160] ,0 ,data[3367:3360] ,data[3375:3368] ,data[3383:3376] ,data[3391:3384] ,0 ,data[3591:3584] ,data[3599:3592] ,data[3607:3600] ,data[3615:3608] ,0 ,data[3815:3808] ,data[3823:3816] ,data[3831:3824] ,data[3839:3832] };
end
422 :begin
 dPIn = {data[2919:2912] ,data[2927:2920] ,data[2935:2928] ,data[2943:2936] ,data[2951:2944] ,data[3143:3136] ,data[3151:3144] ,data[3159:3152] ,data[3167:3160] ,data[3175:3168] ,data[3367:3360] ,data[3375:3368] ,data[3383:3376] ,data[3391:3384] ,data[3399:3392] ,data[3591:3584] ,data[3599:3592] ,data[3607:3600] ,data[3615:3608] ,data[3623:3616] ,data[3815:3808] ,data[3823:3816] ,data[3831:3824] ,data[3839:3832] ,data[3847:3840] };
end
423 :begin
 dPIn = {data[2927:2920] ,data[2935:2928] ,data[2943:2936] ,data[2951:2944] ,data[2959:2952] ,data[3151:3144] ,data[3159:3152] ,data[3167:3160] ,data[3175:3168] ,data[3183:3176] ,data[3375:3368] ,data[3383:3376] ,data[3391:3384] ,data[3399:3392] ,data[3407:3400] ,data[3599:3592] ,data[3607:3600] ,data[3615:3608] ,data[3623:3616] ,data[3631:3624] ,data[3823:3816] ,data[3831:3824] ,data[3839:3832] ,data[3847:3840] ,data[3855:3848] };
end
424 :begin
 dPIn = {data[2935:2928] ,data[2943:2936] ,data[2951:2944] ,data[2959:2952] ,data[2967:2960] ,data[3159:3152] ,data[3167:3160] ,data[3175:3168] ,data[3183:3176] ,data[3191:3184] ,data[3383:3376] ,data[3391:3384] ,data[3399:3392] ,data[3407:3400] ,data[3415:3408] ,data[3607:3600] ,data[3615:3608] ,data[3623:3616] ,data[3631:3624] ,data[3639:3632] ,data[3831:3824] ,data[3839:3832] ,data[3847:3840] ,data[3855:3848] ,data[3863:3856] };
end
425 :begin
 dPIn = {data[2943:2936] ,data[2951:2944] ,data[2959:2952] ,data[2967:2960] ,data[2975:2968] ,data[3167:3160] ,data[3175:3168] ,data[3183:3176] ,data[3191:3184] ,data[3199:3192] ,data[3391:3384] ,data[3399:3392] ,data[3407:3400] ,data[3415:3408] ,data[3423:3416] ,data[3615:3608] ,data[3623:3616] ,data[3631:3624] ,data[3639:3632] ,data[3647:3640] ,data[3839:3832] ,data[3847:3840] ,data[3855:3848] ,data[3863:3856] ,data[3871:3864] };
end
426 :begin
 dPIn = {data[2951:2944] ,data[2959:2952] ,data[2967:2960] ,data[2975:2968] ,data[2983:2976] ,data[3175:3168] ,data[3183:3176] ,data[3191:3184] ,data[3199:3192] ,data[3207:3200] ,data[3399:3392] ,data[3407:3400] ,data[3415:3408] ,data[3423:3416] ,data[3431:3424] ,data[3623:3616] ,data[3631:3624] ,data[3639:3632] ,data[3647:3640] ,data[3655:3648] ,data[3847:3840] ,data[3855:3848] ,data[3863:3856] ,data[3871:3864] ,data[3879:3872] };
end
427 :begin
 dPIn = {data[2959:2952] ,data[2967:2960] ,data[2975:2968] ,data[2983:2976] ,data[2991:2984] ,data[3183:3176] ,data[3191:3184] ,data[3199:3192] ,data[3207:3200] ,data[3215:3208] ,data[3407:3400] ,data[3415:3408] ,data[3423:3416] ,data[3431:3424] ,data[3439:3432] ,data[3631:3624] ,data[3639:3632] ,data[3647:3640] ,data[3655:3648] ,data[3663:3656] ,data[3855:3848] ,data[3863:3856] ,data[3871:3864] ,data[3879:3872] ,data[3887:3880] };
end
428 :begin
 dPIn = {data[2967:2960] ,data[2975:2968] ,data[2983:2976] ,data[2991:2984] ,data[2999:2992] ,data[3191:3184] ,data[3199:3192] ,data[3207:3200] ,data[3215:3208] ,data[3223:3216] ,data[3415:3408] ,data[3423:3416] ,data[3431:3424] ,data[3439:3432] ,data[3447:3440] ,data[3639:3632] ,data[3647:3640] ,data[3655:3648] ,data[3663:3656] ,data[3671:3664] ,data[3863:3856] ,data[3871:3864] ,data[3879:3872] ,data[3887:3880] ,data[3895:3888] };
end
429 :begin
 dPIn = {data[2975:2968] ,data[2983:2976] ,data[2991:2984] ,data[2999:2992] ,data[3007:3000] ,data[3199:3192] ,data[3207:3200] ,data[3215:3208] ,data[3223:3216] ,data[3231:3224] ,data[3423:3416] ,data[3431:3424] ,data[3439:3432] ,data[3447:3440] ,data[3455:3448] ,data[3647:3640] ,data[3655:3648] ,data[3663:3656] ,data[3671:3664] ,data[3679:3672] ,data[3871:3864] ,data[3879:3872] ,data[3887:3880] ,data[3895:3888] ,data[3903:3896] };
end
430 :begin
 dPIn = {data[2983:2976] ,data[2991:2984] ,data[2999:2992] ,data[3007:3000] ,data[3015:3008] ,data[3207:3200] ,data[3215:3208] ,data[3223:3216] ,data[3231:3224] ,data[3239:3232] ,data[3431:3424] ,data[3439:3432] ,data[3447:3440] ,data[3455:3448] ,data[3463:3456] ,data[3655:3648] ,data[3663:3656] ,data[3671:3664] ,data[3679:3672] ,data[3687:3680] ,data[3879:3872] ,data[3887:3880] ,data[3895:3888] ,data[3903:3896] ,data[3911:3904] };
end
431 :begin
 dPIn = {data[2991:2984] ,data[2999:2992] ,data[3007:3000] ,data[3015:3008] ,data[3023:3016] ,data[3215:3208] ,data[3223:3216] ,data[3231:3224] ,data[3239:3232] ,data[3247:3240] ,data[3439:3432] ,data[3447:3440] ,data[3455:3448] ,data[3463:3456] ,data[3471:3464] ,data[3663:3656] ,data[3671:3664] ,data[3679:3672] ,data[3687:3680] ,data[3695:3688] ,data[3887:3880] ,data[3895:3888] ,data[3903:3896] ,data[3911:3904] ,data[3919:3912] };
end
432 :begin
 dPIn = {data[2999:2992] ,data[3007:3000] ,data[3015:3008] ,data[3023:3016] ,data[3031:3024] ,data[3223:3216] ,data[3231:3224] ,data[3239:3232] ,data[3247:3240] ,data[3255:3248] ,data[3447:3440] ,data[3455:3448] ,data[3463:3456] ,data[3471:3464] ,data[3479:3472] ,data[3671:3664] ,data[3679:3672] ,data[3687:3680] ,data[3695:3688] ,data[3703:3696] ,data[3895:3888] ,data[3903:3896] ,data[3911:3904] ,data[3919:3912] ,data[3927:3920] };
end
433 :begin
 dPIn = {data[3007:3000] ,data[3015:3008] ,data[3023:3016] ,data[3031:3024] ,data[3039:3032] ,data[3231:3224] ,data[3239:3232] ,data[3247:3240] ,data[3255:3248] ,data[3263:3256] ,data[3455:3448] ,data[3463:3456] ,data[3471:3464] ,data[3479:3472] ,data[3487:3480] ,data[3679:3672] ,data[3687:3680] ,data[3695:3688] ,data[3703:3696] ,data[3711:3704] ,data[3903:3896] ,data[3911:3904] ,data[3919:3912] ,data[3927:3920] ,data[3935:3928] };
end
434 :begin
 dPIn = {data[3015:3008] ,data[3023:3016] ,data[3031:3024] ,data[3039:3032] ,data[3047:3040] ,data[3239:3232] ,data[3247:3240] ,data[3255:3248] ,data[3263:3256] ,data[3271:3264] ,data[3463:3456] ,data[3471:3464] ,data[3479:3472] ,data[3487:3480] ,data[3495:3488] ,data[3687:3680] ,data[3695:3688] ,data[3703:3696] ,data[3711:3704] ,data[3719:3712] ,data[3911:3904] ,data[3919:3912] ,data[3927:3920] ,data[3935:3928] ,data[3943:3936] };
end
435 :begin
 dPIn = {data[3023:3016] ,data[3031:3024] ,data[3039:3032] ,data[3047:3040] ,data[3055:3048] ,data[3247:3240] ,data[3255:3248] ,data[3263:3256] ,data[3271:3264] ,data[3279:3272] ,data[3471:3464] ,data[3479:3472] ,data[3487:3480] ,data[3495:3488] ,data[3503:3496] ,data[3695:3688] ,data[3703:3696] ,data[3711:3704] ,data[3719:3712] ,data[3727:3720] ,data[3919:3912] ,data[3927:3920] ,data[3935:3928] ,data[3943:3936] ,data[3951:3944] };
end
436 :begin
 dPIn = {data[3031:3024] ,data[3039:3032] ,data[3047:3040] ,data[3055:3048] ,data[3063:3056] ,data[3255:3248] ,data[3263:3256] ,data[3271:3264] ,data[3279:3272] ,data[3287:3280] ,data[3479:3472] ,data[3487:3480] ,data[3495:3488] ,data[3503:3496] ,data[3511:3504] ,data[3703:3696] ,data[3711:3704] ,data[3719:3712] ,data[3727:3720] ,data[3735:3728] ,data[3927:3920] ,data[3935:3928] ,data[3943:3936] ,data[3951:3944] ,data[3959:3952] };
end
437 :begin
 dPIn = {data[3039:3032] ,data[3047:3040] ,data[3055:3048] ,data[3063:3056] ,data[3071:3064] ,data[3263:3256] ,data[3271:3264] ,data[3279:3272] ,data[3287:3280] ,data[3295:3288] ,data[3487:3480] ,data[3495:3488] ,data[3503:3496] ,data[3511:3504] ,data[3519:3512] ,data[3711:3704] ,data[3719:3712] ,data[3727:3720] ,data[3735:3728] ,data[3743:3736] ,data[3935:3928] ,data[3943:3936] ,data[3951:3944] ,data[3959:3952] ,data[3967:3960] };
end
438 :begin
 dPIn = {data[3047:3040] ,data[3055:3048] ,data[3063:3056] ,data[3071:3064] ,data[3079:3072] ,data[3271:3264] ,data[3279:3272] ,data[3287:3280] ,data[3295:3288] ,data[3303:3296] ,data[3495:3488] ,data[3503:3496] ,data[3511:3504] ,data[3519:3512] ,data[3527:3520] ,data[3719:3712] ,data[3727:3720] ,data[3735:3728] ,data[3743:3736] ,data[3751:3744] ,data[3943:3936] ,data[3951:3944] ,data[3959:3952] ,data[3967:3960] ,data[3975:3968] };
end
439 :begin
 dPIn = {data[3055:3048] ,data[3063:3056] ,data[3071:3064] ,data[3079:3072] ,data[3087:3080] ,data[3279:3272] ,data[3287:3280] ,data[3295:3288] ,data[3303:3296] ,data[3311:3304] ,data[3503:3496] ,data[3511:3504] ,data[3519:3512] ,data[3527:3520] ,data[3535:3528] ,data[3727:3720] ,data[3735:3728] ,data[3743:3736] ,data[3751:3744] ,data[3759:3752] ,data[3951:3944] ,data[3959:3952] ,data[3967:3960] ,data[3975:3968] ,data[3983:3976] };
end
440 :begin
 dPIn = {data[3063:3056] ,data[3071:3064] ,data[3079:3072] ,data[3087:3080] ,data[3095:3088] ,data[3287:3280] ,data[3295:3288] ,data[3303:3296] ,data[3311:3304] ,data[3319:3312] ,data[3511:3504] ,data[3519:3512] ,data[3527:3520] ,data[3535:3528] ,data[3543:3536] ,data[3735:3728] ,data[3743:3736] ,data[3751:3744] ,data[3759:3752] ,data[3767:3760] ,data[3959:3952] ,data[3967:3960] ,data[3975:3968] ,data[3983:3976] ,data[3991:3984] };
end
441 :begin
 dPIn = {data[3071:3064] ,data[3079:3072] ,data[3087:3080] ,data[3095:3088] ,data[3103:3096] ,data[3295:3288] ,data[3303:3296] ,data[3311:3304] ,data[3319:3312] ,data[3327:3320] ,data[3519:3512] ,data[3527:3520] ,data[3535:3528] ,data[3543:3536] ,data[3551:3544] ,data[3743:3736] ,data[3751:3744] ,data[3759:3752] ,data[3767:3760] ,data[3775:3768] ,data[3967:3960] ,data[3975:3968] ,data[3983:3976] ,data[3991:3984] ,data[3999:3992] };
end
442 :begin
 dPIn = {data[3079:3072] ,data[3087:3080] ,data[3095:3088] ,data[3103:3096] ,data[3111:3104] ,data[3303:3296] ,data[3311:3304] ,data[3319:3312] ,data[3327:3320] ,data[3335:3328] ,data[3527:3520] ,data[3535:3528] ,data[3543:3536] ,data[3551:3544] ,data[3559:3552] ,data[3751:3744] ,data[3759:3752] ,data[3767:3760] ,data[3775:3768] ,data[3783:3776] ,data[3975:3968] ,data[3983:3976] ,data[3991:3984] ,data[3999:3992] ,data[4007:4000] };
end
443 :begin
 dPIn = {data[3087:3080] ,data[3095:3088] ,data[3103:3096] ,data[3111:3104] ,data[3119:3112] ,data[3311:3304] ,data[3319:3312] ,data[3327:3320] ,data[3335:3328] ,data[3343:3336] ,data[3535:3528] ,data[3543:3536] ,data[3551:3544] ,data[3559:3552] ,data[3567:3560] ,data[3759:3752] ,data[3767:3760] ,data[3775:3768] ,data[3783:3776] ,data[3791:3784] ,data[3983:3976] ,data[3991:3984] ,data[3999:3992] ,data[4007:4000] ,data[4015:4008] };
end
444 :begin
 dPIn = {data[3095:3088] ,data[3103:3096] ,data[3111:3104] ,data[3119:3112] ,data[3127:3120] ,data[3319:3312] ,data[3327:3320] ,data[3335:3328] ,data[3343:3336] ,data[3351:3344] ,data[3543:3536] ,data[3551:3544] ,data[3559:3552] ,data[3567:3560] ,data[3575:3568] ,data[3767:3760] ,data[3775:3768] ,data[3783:3776] ,data[3791:3784] ,data[3799:3792] ,data[3991:3984] ,data[3999:3992] ,data[4007:4000] ,data[4015:4008] ,data[4023:4016] };
end
445 :begin
 dPIn = {data[3103:3096] ,data[3111:3104] ,data[3119:3112] ,data[3127:3120] ,data[3135:3128] ,data[3327:3320] ,data[3335:3328] ,data[3343:3336] ,data[3351:3344] ,data[3359:3352] ,data[3551:3544] ,data[3559:3552] ,data[3567:3560] ,data[3575:3568] ,data[3583:3576] ,data[3775:3768] ,data[3783:3776] ,data[3791:3784] ,data[3799:3792] ,data[3807:3800] ,data[3999:3992] ,data[4007:4000] ,data[4015:4008] ,data[4023:4016] ,data[4031:4024] };
end
446 :begin
 dPIn = {data[3111:3104] ,data[3119:3112] ,data[3127:3120] ,data[3135:3128] ,0 ,data[3335:3328] ,data[3343:3336] ,data[3351:3344] ,data[3359:3352] ,0 ,data[3559:3552] ,data[3567:3560] ,data[3575:3568] ,data[3583:3576] ,0 ,data[3783:3776] ,data[3791:3784] ,data[3799:3792] ,data[3807:3800] ,0 ,data[4007:4000] ,data[4015:4008] ,data[4023:4016] ,data[4031:4024] ,0 };
end
447 :begin
 dPIn = {data[3119:3112] ,data[3127:3120] ,data[3135:3128] ,0 ,0 ,data[3343:3336] ,data[3351:3344] ,data[3359:3352] ,0 ,0 ,data[3567:3560] ,data[3575:3568] ,data[3583:3576] ,0 ,0 ,data[3791:3784] ,data[3799:3792] ,data[3807:3800] ,0 ,0 ,data[4015:4008] ,data[4023:4016] ,data[4031:4024] ,0 ,0 };
end
448 :begin
 dPIn = {0 ,0 ,data[3143:3136] ,data[3151:3144] ,data[3159:3152] ,0 ,0 ,data[3367:3360] ,data[3375:3368] ,data[3383:3376] ,0 ,0 ,data[3591:3584] ,data[3599:3592] ,data[3607:3600] ,0 ,0 ,data[3815:3808] ,data[3823:3816] ,data[3831:3824] ,0 ,0 ,data[4039:4032] ,data[4047:4040] ,data[4055:4048] };
end
449 :begin
 dPIn = {0 ,data[3143:3136] ,data[3151:3144] ,data[3159:3152] ,data[3167:3160] ,0 ,data[3367:3360] ,data[3375:3368] ,data[3383:3376] ,data[3391:3384] ,0 ,data[3591:3584] ,data[3599:3592] ,data[3607:3600] ,data[3615:3608] ,0 ,data[3815:3808] ,data[3823:3816] ,data[3831:3824] ,data[3839:3832] ,0 ,data[4039:4032] ,data[4047:4040] ,data[4055:4048] ,data[4063:4056] };
end
450 :begin
 dPIn = {data[3143:3136] ,data[3151:3144] ,data[3159:3152] ,data[3167:3160] ,data[3175:3168] ,data[3367:3360] ,data[3375:3368] ,data[3383:3376] ,data[3391:3384] ,data[3399:3392] ,data[3591:3584] ,data[3599:3592] ,data[3607:3600] ,data[3615:3608] ,data[3623:3616] ,data[3815:3808] ,data[3823:3816] ,data[3831:3824] ,data[3839:3832] ,data[3847:3840] ,data[4039:4032] ,data[4047:4040] ,data[4055:4048] ,data[4063:4056] ,data[4071:4064] };
end
451 :begin
 dPIn = {data[3151:3144] ,data[3159:3152] ,data[3167:3160] ,data[3175:3168] ,data[3183:3176] ,data[3375:3368] ,data[3383:3376] ,data[3391:3384] ,data[3399:3392] ,data[3407:3400] ,data[3599:3592] ,data[3607:3600] ,data[3615:3608] ,data[3623:3616] ,data[3631:3624] ,data[3823:3816] ,data[3831:3824] ,data[3839:3832] ,data[3847:3840] ,data[3855:3848] ,data[4047:4040] ,data[4055:4048] ,data[4063:4056] ,data[4071:4064] ,data[4079:4072] };
end
452 :begin
 dPIn = {data[3159:3152] ,data[3167:3160] ,data[3175:3168] ,data[3183:3176] ,data[3191:3184] ,data[3383:3376] ,data[3391:3384] ,data[3399:3392] ,data[3407:3400] ,data[3415:3408] ,data[3607:3600] ,data[3615:3608] ,data[3623:3616] ,data[3631:3624] ,data[3639:3632] ,data[3831:3824] ,data[3839:3832] ,data[3847:3840] ,data[3855:3848] ,data[3863:3856] ,data[4055:4048] ,data[4063:4056] ,data[4071:4064] ,data[4079:4072] ,data[4087:4080] };
end
453 :begin
 dPIn = {data[3167:3160] ,data[3175:3168] ,data[3183:3176] ,data[3191:3184] ,data[3199:3192] ,data[3391:3384] ,data[3399:3392] ,data[3407:3400] ,data[3415:3408] ,data[3423:3416] ,data[3615:3608] ,data[3623:3616] ,data[3631:3624] ,data[3639:3632] ,data[3647:3640] ,data[3839:3832] ,data[3847:3840] ,data[3855:3848] ,data[3863:3856] ,data[3871:3864] ,data[4063:4056] ,data[4071:4064] ,data[4079:4072] ,data[4087:4080] ,data[4095:4088] };
end
454 :begin
 dPIn = {data[3175:3168] ,data[3183:3176] ,data[3191:3184] ,data[3199:3192] ,data[3207:3200] ,data[3399:3392] ,data[3407:3400] ,data[3415:3408] ,data[3423:3416] ,data[3431:3424] ,data[3623:3616] ,data[3631:3624] ,data[3639:3632] ,data[3647:3640] ,data[3655:3648] ,data[3847:3840] ,data[3855:3848] ,data[3863:3856] ,data[3871:3864] ,data[3879:3872] ,data[4071:4064] ,data[4079:4072] ,data[4087:4080] ,data[4095:4088] ,data[4103:4096] };
end
455 :begin
 dPIn = {data[3183:3176] ,data[3191:3184] ,data[3199:3192] ,data[3207:3200] ,data[3215:3208] ,data[3407:3400] ,data[3415:3408] ,data[3423:3416] ,data[3431:3424] ,data[3439:3432] ,data[3631:3624] ,data[3639:3632] ,data[3647:3640] ,data[3655:3648] ,data[3663:3656] ,data[3855:3848] ,data[3863:3856] ,data[3871:3864] ,data[3879:3872] ,data[3887:3880] ,data[4079:4072] ,data[4087:4080] ,data[4095:4088] ,data[4103:4096] ,data[4111:4104] };
end
456 :begin
 dPIn = {data[3191:3184] ,data[3199:3192] ,data[3207:3200] ,data[3215:3208] ,data[3223:3216] ,data[3415:3408] ,data[3423:3416] ,data[3431:3424] ,data[3439:3432] ,data[3447:3440] ,data[3639:3632] ,data[3647:3640] ,data[3655:3648] ,data[3663:3656] ,data[3671:3664] ,data[3863:3856] ,data[3871:3864] ,data[3879:3872] ,data[3887:3880] ,data[3895:3888] ,data[4087:4080] ,data[4095:4088] ,data[4103:4096] ,data[4111:4104] ,data[4119:4112] };
end
457 :begin
 dPIn = {data[3199:3192] ,data[3207:3200] ,data[3215:3208] ,data[3223:3216] ,data[3231:3224] ,data[3423:3416] ,data[3431:3424] ,data[3439:3432] ,data[3447:3440] ,data[3455:3448] ,data[3647:3640] ,data[3655:3648] ,data[3663:3656] ,data[3671:3664] ,data[3679:3672] ,data[3871:3864] ,data[3879:3872] ,data[3887:3880] ,data[3895:3888] ,data[3903:3896] ,data[4095:4088] ,data[4103:4096] ,data[4111:4104] ,data[4119:4112] ,data[4127:4120] };
end
458 :begin
 dPIn = {data[3207:3200] ,data[3215:3208] ,data[3223:3216] ,data[3231:3224] ,data[3239:3232] ,data[3431:3424] ,data[3439:3432] ,data[3447:3440] ,data[3455:3448] ,data[3463:3456] ,data[3655:3648] ,data[3663:3656] ,data[3671:3664] ,data[3679:3672] ,data[3687:3680] ,data[3879:3872] ,data[3887:3880] ,data[3895:3888] ,data[3903:3896] ,data[3911:3904] ,data[4103:4096] ,data[4111:4104] ,data[4119:4112] ,data[4127:4120] ,data[4135:4128] };
end
459 :begin
 dPIn = {data[3215:3208] ,data[3223:3216] ,data[3231:3224] ,data[3239:3232] ,data[3247:3240] ,data[3439:3432] ,data[3447:3440] ,data[3455:3448] ,data[3463:3456] ,data[3471:3464] ,data[3663:3656] ,data[3671:3664] ,data[3679:3672] ,data[3687:3680] ,data[3695:3688] ,data[3887:3880] ,data[3895:3888] ,data[3903:3896] ,data[3911:3904] ,data[3919:3912] ,data[4111:4104] ,data[4119:4112] ,data[4127:4120] ,data[4135:4128] ,data[4143:4136] };
end
460 :begin
 dPIn = {data[3223:3216] ,data[3231:3224] ,data[3239:3232] ,data[3247:3240] ,data[3255:3248] ,data[3447:3440] ,data[3455:3448] ,data[3463:3456] ,data[3471:3464] ,data[3479:3472] ,data[3671:3664] ,data[3679:3672] ,data[3687:3680] ,data[3695:3688] ,data[3703:3696] ,data[3895:3888] ,data[3903:3896] ,data[3911:3904] ,data[3919:3912] ,data[3927:3920] ,data[4119:4112] ,data[4127:4120] ,data[4135:4128] ,data[4143:4136] ,data[4151:4144] };
end
461 :begin
 dPIn = {data[3231:3224] ,data[3239:3232] ,data[3247:3240] ,data[3255:3248] ,data[3263:3256] ,data[3455:3448] ,data[3463:3456] ,data[3471:3464] ,data[3479:3472] ,data[3487:3480] ,data[3679:3672] ,data[3687:3680] ,data[3695:3688] ,data[3703:3696] ,data[3711:3704] ,data[3903:3896] ,data[3911:3904] ,data[3919:3912] ,data[3927:3920] ,data[3935:3928] ,data[4127:4120] ,data[4135:4128] ,data[4143:4136] ,data[4151:4144] ,data[4159:4152] };
end
462 :begin
 dPIn = {data[3239:3232] ,data[3247:3240] ,data[3255:3248] ,data[3263:3256] ,data[3271:3264] ,data[3463:3456] ,data[3471:3464] ,data[3479:3472] ,data[3487:3480] ,data[3495:3488] ,data[3687:3680] ,data[3695:3688] ,data[3703:3696] ,data[3711:3704] ,data[3719:3712] ,data[3911:3904] ,data[3919:3912] ,data[3927:3920] ,data[3935:3928] ,data[3943:3936] ,data[4135:4128] ,data[4143:4136] ,data[4151:4144] ,data[4159:4152] ,data[4167:4160] };
end
463 :begin
 dPIn = {data[3247:3240] ,data[3255:3248] ,data[3263:3256] ,data[3271:3264] ,data[3279:3272] ,data[3471:3464] ,data[3479:3472] ,data[3487:3480] ,data[3495:3488] ,data[3503:3496] ,data[3695:3688] ,data[3703:3696] ,data[3711:3704] ,data[3719:3712] ,data[3727:3720] ,data[3919:3912] ,data[3927:3920] ,data[3935:3928] ,data[3943:3936] ,data[3951:3944] ,data[4143:4136] ,data[4151:4144] ,data[4159:4152] ,data[4167:4160] ,data[4175:4168] };
end
464 :begin
 dPIn = {data[3255:3248] ,data[3263:3256] ,data[3271:3264] ,data[3279:3272] ,data[3287:3280] ,data[3479:3472] ,data[3487:3480] ,data[3495:3488] ,data[3503:3496] ,data[3511:3504] ,data[3703:3696] ,data[3711:3704] ,data[3719:3712] ,data[3727:3720] ,data[3735:3728] ,data[3927:3920] ,data[3935:3928] ,data[3943:3936] ,data[3951:3944] ,data[3959:3952] ,data[4151:4144] ,data[4159:4152] ,data[4167:4160] ,data[4175:4168] ,data[4183:4176] };
end
465 :begin
 dPIn = {data[3263:3256] ,data[3271:3264] ,data[3279:3272] ,data[3287:3280] ,data[3295:3288] ,data[3487:3480] ,data[3495:3488] ,data[3503:3496] ,data[3511:3504] ,data[3519:3512] ,data[3711:3704] ,data[3719:3712] ,data[3727:3720] ,data[3735:3728] ,data[3743:3736] ,data[3935:3928] ,data[3943:3936] ,data[3951:3944] ,data[3959:3952] ,data[3967:3960] ,data[4159:4152] ,data[4167:4160] ,data[4175:4168] ,data[4183:4176] ,data[4191:4184] };
end
466 :begin
 dPIn = {data[3271:3264] ,data[3279:3272] ,data[3287:3280] ,data[3295:3288] ,data[3303:3296] ,data[3495:3488] ,data[3503:3496] ,data[3511:3504] ,data[3519:3512] ,data[3527:3520] ,data[3719:3712] ,data[3727:3720] ,data[3735:3728] ,data[3743:3736] ,data[3751:3744] ,data[3943:3936] ,data[3951:3944] ,data[3959:3952] ,data[3967:3960] ,data[3975:3968] ,data[4167:4160] ,data[4175:4168] ,data[4183:4176] ,data[4191:4184] ,data[4199:4192] };
end
467 :begin
 dPIn = {data[3279:3272] ,data[3287:3280] ,data[3295:3288] ,data[3303:3296] ,data[3311:3304] ,data[3503:3496] ,data[3511:3504] ,data[3519:3512] ,data[3527:3520] ,data[3535:3528] ,data[3727:3720] ,data[3735:3728] ,data[3743:3736] ,data[3751:3744] ,data[3759:3752] ,data[3951:3944] ,data[3959:3952] ,data[3967:3960] ,data[3975:3968] ,data[3983:3976] ,data[4175:4168] ,data[4183:4176] ,data[4191:4184] ,data[4199:4192] ,data[4207:4200] };
end
468 :begin
 dPIn = {data[3287:3280] ,data[3295:3288] ,data[3303:3296] ,data[3311:3304] ,data[3319:3312] ,data[3511:3504] ,data[3519:3512] ,data[3527:3520] ,data[3535:3528] ,data[3543:3536] ,data[3735:3728] ,data[3743:3736] ,data[3751:3744] ,data[3759:3752] ,data[3767:3760] ,data[3959:3952] ,data[3967:3960] ,data[3975:3968] ,data[3983:3976] ,data[3991:3984] ,data[4183:4176] ,data[4191:4184] ,data[4199:4192] ,data[4207:4200] ,data[4215:4208] };
end
469 :begin
 dPIn = {data[3295:3288] ,data[3303:3296] ,data[3311:3304] ,data[3319:3312] ,data[3327:3320] ,data[3519:3512] ,data[3527:3520] ,data[3535:3528] ,data[3543:3536] ,data[3551:3544] ,data[3743:3736] ,data[3751:3744] ,data[3759:3752] ,data[3767:3760] ,data[3775:3768] ,data[3967:3960] ,data[3975:3968] ,data[3983:3976] ,data[3991:3984] ,data[3999:3992] ,data[4191:4184] ,data[4199:4192] ,data[4207:4200] ,data[4215:4208] ,data[4223:4216] };
end
470 :begin
 dPIn = {data[3303:3296] ,data[3311:3304] ,data[3319:3312] ,data[3327:3320] ,data[3335:3328] ,data[3527:3520] ,data[3535:3528] ,data[3543:3536] ,data[3551:3544] ,data[3559:3552] ,data[3751:3744] ,data[3759:3752] ,data[3767:3760] ,data[3775:3768] ,data[3783:3776] ,data[3975:3968] ,data[3983:3976] ,data[3991:3984] ,data[3999:3992] ,data[4007:4000] ,data[4199:4192] ,data[4207:4200] ,data[4215:4208] ,data[4223:4216] ,data[4231:4224] };
end
471 :begin
 dPIn = {data[3311:3304] ,data[3319:3312] ,data[3327:3320] ,data[3335:3328] ,data[3343:3336] ,data[3535:3528] ,data[3543:3536] ,data[3551:3544] ,data[3559:3552] ,data[3567:3560] ,data[3759:3752] ,data[3767:3760] ,data[3775:3768] ,data[3783:3776] ,data[3791:3784] ,data[3983:3976] ,data[3991:3984] ,data[3999:3992] ,data[4007:4000] ,data[4015:4008] ,data[4207:4200] ,data[4215:4208] ,data[4223:4216] ,data[4231:4224] ,data[4239:4232] };
end
472 :begin
 dPIn = {data[3319:3312] ,data[3327:3320] ,data[3335:3328] ,data[3343:3336] ,data[3351:3344] ,data[3543:3536] ,data[3551:3544] ,data[3559:3552] ,data[3567:3560] ,data[3575:3568] ,data[3767:3760] ,data[3775:3768] ,data[3783:3776] ,data[3791:3784] ,data[3799:3792] ,data[3991:3984] ,data[3999:3992] ,data[4007:4000] ,data[4015:4008] ,data[4023:4016] ,data[4215:4208] ,data[4223:4216] ,data[4231:4224] ,data[4239:4232] ,data[4247:4240] };
end
473 :begin
 dPIn = {data[3327:3320] ,data[3335:3328] ,data[3343:3336] ,data[3351:3344] ,data[3359:3352] ,data[3551:3544] ,data[3559:3552] ,data[3567:3560] ,data[3575:3568] ,data[3583:3576] ,data[3775:3768] ,data[3783:3776] ,data[3791:3784] ,data[3799:3792] ,data[3807:3800] ,data[3999:3992] ,data[4007:4000] ,data[4015:4008] ,data[4023:4016] ,data[4031:4024] ,data[4223:4216] ,data[4231:4224] ,data[4239:4232] ,data[4247:4240] ,data[4255:4248] };
end
474 :begin
 dPIn = {data[3335:3328] ,data[3343:3336] ,data[3351:3344] ,data[3359:3352] ,0 ,data[3559:3552] ,data[3567:3560] ,data[3575:3568] ,data[3583:3576] ,0 ,data[3783:3776] ,data[3791:3784] ,data[3799:3792] ,data[3807:3800] ,0 ,data[4007:4000] ,data[4015:4008] ,data[4023:4016] ,data[4031:4024] ,0 ,data[4231:4224] ,data[4239:4232] ,data[4247:4240] ,data[4255:4248] ,0 };
end
475 :begin
 dPIn = {data[3343:3336] ,data[3351:3344] ,data[3359:3352] ,0 ,0 ,data[3567:3560] ,data[3575:3568] ,data[3583:3576] ,0 ,0 ,data[3791:3784] ,data[3799:3792] ,data[3807:3800] ,0 ,0 ,data[4015:4008] ,data[4023:4016] ,data[4031:4024] ,0 ,0 ,data[4239:4232] ,data[4247:4240] ,data[4255:4248] ,0 ,0 };
end
476 :begin
 dPIn = {0 ,0 ,data[3367:3360] ,data[3375:3368] ,data[3383:3376] ,0 ,0 ,data[3591:3584] ,data[3599:3592] ,data[3607:3600] ,0 ,0 ,data[3815:3808] ,data[3823:3816] ,data[3831:3824] ,0 ,0 ,data[4039:4032] ,data[4047:4040] ,data[4055:4048] ,0 ,0 ,data[4263:4256] ,data[4271:4264] ,data[4279:4272] };
end
477 :begin
 dPIn = {0 ,data[3367:3360] ,data[3375:3368] ,data[3383:3376] ,data[3391:3384] ,0 ,data[3591:3584] ,data[3599:3592] ,data[3607:3600] ,data[3615:3608] ,0 ,data[3815:3808] ,data[3823:3816] ,data[3831:3824] ,data[3839:3832] ,0 ,data[4039:4032] ,data[4047:4040] ,data[4055:4048] ,data[4063:4056] ,0 ,data[4263:4256] ,data[4271:4264] ,data[4279:4272] ,data[4287:4280] };
end
478 :begin
 dPIn = {data[3367:3360] ,data[3375:3368] ,data[3383:3376] ,data[3391:3384] ,data[3399:3392] ,data[3591:3584] ,data[3599:3592] ,data[3607:3600] ,data[3615:3608] ,data[3623:3616] ,data[3815:3808] ,data[3823:3816] ,data[3831:3824] ,data[3839:3832] ,data[3847:3840] ,data[4039:4032] ,data[4047:4040] ,data[4055:4048] ,data[4063:4056] ,data[4071:4064] ,data[4263:4256] ,data[4271:4264] ,data[4279:4272] ,data[4287:4280] ,data[4295:4288] };
end
479 :begin
 dPIn = {data[3375:3368] ,data[3383:3376] ,data[3391:3384] ,data[3399:3392] ,data[3407:3400] ,data[3599:3592] ,data[3607:3600] ,data[3615:3608] ,data[3623:3616] ,data[3631:3624] ,data[3823:3816] ,data[3831:3824] ,data[3839:3832] ,data[3847:3840] ,data[3855:3848] ,data[4047:4040] ,data[4055:4048] ,data[4063:4056] ,data[4071:4064] ,data[4079:4072] ,data[4271:4264] ,data[4279:4272] ,data[4287:4280] ,data[4295:4288] ,data[4303:4296] };
end
480 :begin
 dPIn = {data[3383:3376] ,data[3391:3384] ,data[3399:3392] ,data[3407:3400] ,data[3415:3408] ,data[3607:3600] ,data[3615:3608] ,data[3623:3616] ,data[3631:3624] ,data[3639:3632] ,data[3831:3824] ,data[3839:3832] ,data[3847:3840] ,data[3855:3848] ,data[3863:3856] ,data[4055:4048] ,data[4063:4056] ,data[4071:4064] ,data[4079:4072] ,data[4087:4080] ,data[4279:4272] ,data[4287:4280] ,data[4295:4288] ,data[4303:4296] ,data[4311:4304] };
end
481 :begin
 dPIn = {data[3391:3384] ,data[3399:3392] ,data[3407:3400] ,data[3415:3408] ,data[3423:3416] ,data[3615:3608] ,data[3623:3616] ,data[3631:3624] ,data[3639:3632] ,data[3647:3640] ,data[3839:3832] ,data[3847:3840] ,data[3855:3848] ,data[3863:3856] ,data[3871:3864] ,data[4063:4056] ,data[4071:4064] ,data[4079:4072] ,data[4087:4080] ,data[4095:4088] ,data[4287:4280] ,data[4295:4288] ,data[4303:4296] ,data[4311:4304] ,data[4319:4312] };
end
482 :begin
 dPIn = {data[3399:3392] ,data[3407:3400] ,data[3415:3408] ,data[3423:3416] ,data[3431:3424] ,data[3623:3616] ,data[3631:3624] ,data[3639:3632] ,data[3647:3640] ,data[3655:3648] ,data[3847:3840] ,data[3855:3848] ,data[3863:3856] ,data[3871:3864] ,data[3879:3872] ,data[4071:4064] ,data[4079:4072] ,data[4087:4080] ,data[4095:4088] ,data[4103:4096] ,data[4295:4288] ,data[4303:4296] ,data[4311:4304] ,data[4319:4312] ,data[4327:4320] };
end
483 :begin
 dPIn = {data[3407:3400] ,data[3415:3408] ,data[3423:3416] ,data[3431:3424] ,data[3439:3432] ,data[3631:3624] ,data[3639:3632] ,data[3647:3640] ,data[3655:3648] ,data[3663:3656] ,data[3855:3848] ,data[3863:3856] ,data[3871:3864] ,data[3879:3872] ,data[3887:3880] ,data[4079:4072] ,data[4087:4080] ,data[4095:4088] ,data[4103:4096] ,data[4111:4104] ,data[4303:4296] ,data[4311:4304] ,data[4319:4312] ,data[4327:4320] ,data[4335:4328] };
end
484 :begin
 dPIn = {data[3415:3408] ,data[3423:3416] ,data[3431:3424] ,data[3439:3432] ,data[3447:3440] ,data[3639:3632] ,data[3647:3640] ,data[3655:3648] ,data[3663:3656] ,data[3671:3664] ,data[3863:3856] ,data[3871:3864] ,data[3879:3872] ,data[3887:3880] ,data[3895:3888] ,data[4087:4080] ,data[4095:4088] ,data[4103:4096] ,data[4111:4104] ,data[4119:4112] ,data[4311:4304] ,data[4319:4312] ,data[4327:4320] ,data[4335:4328] ,data[4343:4336] };
end
485 :begin
 dPIn = {data[3423:3416] ,data[3431:3424] ,data[3439:3432] ,data[3447:3440] ,data[3455:3448] ,data[3647:3640] ,data[3655:3648] ,data[3663:3656] ,data[3671:3664] ,data[3679:3672] ,data[3871:3864] ,data[3879:3872] ,data[3887:3880] ,data[3895:3888] ,data[3903:3896] ,data[4095:4088] ,data[4103:4096] ,data[4111:4104] ,data[4119:4112] ,data[4127:4120] ,data[4319:4312] ,data[4327:4320] ,data[4335:4328] ,data[4343:4336] ,data[4351:4344] };
end
486 :begin
 dPIn = {data[3431:3424] ,data[3439:3432] ,data[3447:3440] ,data[3455:3448] ,data[3463:3456] ,data[3655:3648] ,data[3663:3656] ,data[3671:3664] ,data[3679:3672] ,data[3687:3680] ,data[3879:3872] ,data[3887:3880] ,data[3895:3888] ,data[3903:3896] ,data[3911:3904] ,data[4103:4096] ,data[4111:4104] ,data[4119:4112] ,data[4127:4120] ,data[4135:4128] ,data[4327:4320] ,data[4335:4328] ,data[4343:4336] ,data[4351:4344] ,data[4359:4352] };
end
487 :begin
 dPIn = {data[3439:3432] ,data[3447:3440] ,data[3455:3448] ,data[3463:3456] ,data[3471:3464] ,data[3663:3656] ,data[3671:3664] ,data[3679:3672] ,data[3687:3680] ,data[3695:3688] ,data[3887:3880] ,data[3895:3888] ,data[3903:3896] ,data[3911:3904] ,data[3919:3912] ,data[4111:4104] ,data[4119:4112] ,data[4127:4120] ,data[4135:4128] ,data[4143:4136] ,data[4335:4328] ,data[4343:4336] ,data[4351:4344] ,data[4359:4352] ,data[4367:4360] };
end
488 :begin
 dPIn = {data[3447:3440] ,data[3455:3448] ,data[3463:3456] ,data[3471:3464] ,data[3479:3472] ,data[3671:3664] ,data[3679:3672] ,data[3687:3680] ,data[3695:3688] ,data[3703:3696] ,data[3895:3888] ,data[3903:3896] ,data[3911:3904] ,data[3919:3912] ,data[3927:3920] ,data[4119:4112] ,data[4127:4120] ,data[4135:4128] ,data[4143:4136] ,data[4151:4144] ,data[4343:4336] ,data[4351:4344] ,data[4359:4352] ,data[4367:4360] ,data[4375:4368] };
end
489 :begin
 dPIn = {data[3455:3448] ,data[3463:3456] ,data[3471:3464] ,data[3479:3472] ,data[3487:3480] ,data[3679:3672] ,data[3687:3680] ,data[3695:3688] ,data[3703:3696] ,data[3711:3704] ,data[3903:3896] ,data[3911:3904] ,data[3919:3912] ,data[3927:3920] ,data[3935:3928] ,data[4127:4120] ,data[4135:4128] ,data[4143:4136] ,data[4151:4144] ,data[4159:4152] ,data[4351:4344] ,data[4359:4352] ,data[4367:4360] ,data[4375:4368] ,data[4383:4376] };
end
490 :begin
 dPIn = {data[3463:3456] ,data[3471:3464] ,data[3479:3472] ,data[3487:3480] ,data[3495:3488] ,data[3687:3680] ,data[3695:3688] ,data[3703:3696] ,data[3711:3704] ,data[3719:3712] ,data[3911:3904] ,data[3919:3912] ,data[3927:3920] ,data[3935:3928] ,data[3943:3936] ,data[4135:4128] ,data[4143:4136] ,data[4151:4144] ,data[4159:4152] ,data[4167:4160] ,data[4359:4352] ,data[4367:4360] ,data[4375:4368] ,data[4383:4376] ,data[4391:4384] };
end
491 :begin
 dPIn = {data[3471:3464] ,data[3479:3472] ,data[3487:3480] ,data[3495:3488] ,data[3503:3496] ,data[3695:3688] ,data[3703:3696] ,data[3711:3704] ,data[3719:3712] ,data[3727:3720] ,data[3919:3912] ,data[3927:3920] ,data[3935:3928] ,data[3943:3936] ,data[3951:3944] ,data[4143:4136] ,data[4151:4144] ,data[4159:4152] ,data[4167:4160] ,data[4175:4168] ,data[4367:4360] ,data[4375:4368] ,data[4383:4376] ,data[4391:4384] ,data[4399:4392] };
end
492 :begin
 dPIn = {data[3479:3472] ,data[3487:3480] ,data[3495:3488] ,data[3503:3496] ,data[3511:3504] ,data[3703:3696] ,data[3711:3704] ,data[3719:3712] ,data[3727:3720] ,data[3735:3728] ,data[3927:3920] ,data[3935:3928] ,data[3943:3936] ,data[3951:3944] ,data[3959:3952] ,data[4151:4144] ,data[4159:4152] ,data[4167:4160] ,data[4175:4168] ,data[4183:4176] ,data[4375:4368] ,data[4383:4376] ,data[4391:4384] ,data[4399:4392] ,data[4407:4400] };
end
493 :begin
 dPIn = {data[3487:3480] ,data[3495:3488] ,data[3503:3496] ,data[3511:3504] ,data[3519:3512] ,data[3711:3704] ,data[3719:3712] ,data[3727:3720] ,data[3735:3728] ,data[3743:3736] ,data[3935:3928] ,data[3943:3936] ,data[3951:3944] ,data[3959:3952] ,data[3967:3960] ,data[4159:4152] ,data[4167:4160] ,data[4175:4168] ,data[4183:4176] ,data[4191:4184] ,data[4383:4376] ,data[4391:4384] ,data[4399:4392] ,data[4407:4400] ,data[4415:4408] };
end
494 :begin
 dPIn = {data[3495:3488] ,data[3503:3496] ,data[3511:3504] ,data[3519:3512] ,data[3527:3520] ,data[3719:3712] ,data[3727:3720] ,data[3735:3728] ,data[3743:3736] ,data[3751:3744] ,data[3943:3936] ,data[3951:3944] ,data[3959:3952] ,data[3967:3960] ,data[3975:3968] ,data[4167:4160] ,data[4175:4168] ,data[4183:4176] ,data[4191:4184] ,data[4199:4192] ,data[4391:4384] ,data[4399:4392] ,data[4407:4400] ,data[4415:4408] ,data[4423:4416] };
end
495 :begin
 dPIn = {data[3503:3496] ,data[3511:3504] ,data[3519:3512] ,data[3527:3520] ,data[3535:3528] ,data[3727:3720] ,data[3735:3728] ,data[3743:3736] ,data[3751:3744] ,data[3759:3752] ,data[3951:3944] ,data[3959:3952] ,data[3967:3960] ,data[3975:3968] ,data[3983:3976] ,data[4175:4168] ,data[4183:4176] ,data[4191:4184] ,data[4199:4192] ,data[4207:4200] ,data[4399:4392] ,data[4407:4400] ,data[4415:4408] ,data[4423:4416] ,data[4431:4424] };
end
496 :begin
 dPIn = {data[3511:3504] ,data[3519:3512] ,data[3527:3520] ,data[3535:3528] ,data[3543:3536] ,data[3735:3728] ,data[3743:3736] ,data[3751:3744] ,data[3759:3752] ,data[3767:3760] ,data[3959:3952] ,data[3967:3960] ,data[3975:3968] ,data[3983:3976] ,data[3991:3984] ,data[4183:4176] ,data[4191:4184] ,data[4199:4192] ,data[4207:4200] ,data[4215:4208] ,data[4407:4400] ,data[4415:4408] ,data[4423:4416] ,data[4431:4424] ,data[4439:4432] };
end
497 :begin
 dPIn = {data[3519:3512] ,data[3527:3520] ,data[3535:3528] ,data[3543:3536] ,data[3551:3544] ,data[3743:3736] ,data[3751:3744] ,data[3759:3752] ,data[3767:3760] ,data[3775:3768] ,data[3967:3960] ,data[3975:3968] ,data[3983:3976] ,data[3991:3984] ,data[3999:3992] ,data[4191:4184] ,data[4199:4192] ,data[4207:4200] ,data[4215:4208] ,data[4223:4216] ,data[4415:4408] ,data[4423:4416] ,data[4431:4424] ,data[4439:4432] ,data[4447:4440] };
end
498 :begin
 dPIn = {data[3527:3520] ,data[3535:3528] ,data[3543:3536] ,data[3551:3544] ,data[3559:3552] ,data[3751:3744] ,data[3759:3752] ,data[3767:3760] ,data[3775:3768] ,data[3783:3776] ,data[3975:3968] ,data[3983:3976] ,data[3991:3984] ,data[3999:3992] ,data[4007:4000] ,data[4199:4192] ,data[4207:4200] ,data[4215:4208] ,data[4223:4216] ,data[4231:4224] ,data[4423:4416] ,data[4431:4424] ,data[4439:4432] ,data[4447:4440] ,data[4455:4448] };
end
499 :begin
 dPIn = {data[3535:3528] ,data[3543:3536] ,data[3551:3544] ,data[3559:3552] ,data[3567:3560] ,data[3759:3752] ,data[3767:3760] ,data[3775:3768] ,data[3783:3776] ,data[3791:3784] ,data[3983:3976] ,data[3991:3984] ,data[3999:3992] ,data[4007:4000] ,data[4015:4008] ,data[4207:4200] ,data[4215:4208] ,data[4223:4216] ,data[4231:4224] ,data[4239:4232] ,data[4431:4424] ,data[4439:4432] ,data[4447:4440] ,data[4455:4448] ,data[4463:4456] };
end
500 :begin
 dPIn = {data[3543:3536] ,data[3551:3544] ,data[3559:3552] ,data[3567:3560] ,data[3575:3568] ,data[3767:3760] ,data[3775:3768] ,data[3783:3776] ,data[3791:3784] ,data[3799:3792] ,data[3991:3984] ,data[3999:3992] ,data[4007:4000] ,data[4015:4008] ,data[4023:4016] ,data[4215:4208] ,data[4223:4216] ,data[4231:4224] ,data[4239:4232] ,data[4247:4240] ,data[4439:4432] ,data[4447:4440] ,data[4455:4448] ,data[4463:4456] ,data[4471:4464] };
end
501 :begin
 dPIn = {data[3551:3544] ,data[3559:3552] ,data[3567:3560] ,data[3575:3568] ,data[3583:3576] ,data[3775:3768] ,data[3783:3776] ,data[3791:3784] ,data[3799:3792] ,data[3807:3800] ,data[3999:3992] ,data[4007:4000] ,data[4015:4008] ,data[4023:4016] ,data[4031:4024] ,data[4223:4216] ,data[4231:4224] ,data[4239:4232] ,data[4247:4240] ,data[4255:4248] ,data[4447:4440] ,data[4455:4448] ,data[4463:4456] ,data[4471:4464] ,data[4479:4472] };
end
502 :begin
 dPIn = {data[3559:3552] ,data[3567:3560] ,data[3575:3568] ,data[3583:3576] ,0 ,data[3783:3776] ,data[3791:3784] ,data[3799:3792] ,data[3807:3800] ,0 ,data[4007:4000] ,data[4015:4008] ,data[4023:4016] ,data[4031:4024] ,0 ,data[4231:4224] ,data[4239:4232] ,data[4247:4240] ,data[4255:4248] ,0 ,data[4455:4448] ,data[4463:4456] ,data[4471:4464] ,data[4479:4472] ,0 };
end
503 :begin
 dPIn = {data[3567:3560] ,data[3575:3568] ,data[3583:3576] ,0 ,0 ,data[3791:3784] ,data[3799:3792] ,data[3807:3800] ,0 ,0 ,data[4015:4008] ,data[4023:4016] ,data[4031:4024] ,0 ,0 ,data[4239:4232] ,data[4247:4240] ,data[4255:4248] ,0 ,0 ,data[4463:4456] ,data[4471:4464] ,data[4479:4472] ,0 ,0 };
end
504 :begin
 dPIn = {0 ,0 ,data[3591:3584] ,data[3599:3592] ,data[3607:3600] ,0 ,0 ,data[3815:3808] ,data[3823:3816] ,data[3831:3824] ,0 ,0 ,data[4039:4032] ,data[4047:4040] ,data[4055:4048] ,0 ,0 ,data[4263:4256] ,data[4271:4264] ,data[4279:4272] ,0 ,0 ,data[4487:4480] ,data[4495:4488] ,data[4503:4496] };
end
505 :begin
 dPIn = {0 ,data[3591:3584] ,data[3599:3592] ,data[3607:3600] ,data[3615:3608] ,0 ,data[3815:3808] ,data[3823:3816] ,data[3831:3824] ,data[3839:3832] ,0 ,data[4039:4032] ,data[4047:4040] ,data[4055:4048] ,data[4063:4056] ,0 ,data[4263:4256] ,data[4271:4264] ,data[4279:4272] ,data[4287:4280] ,0 ,data[4487:4480] ,data[4495:4488] ,data[4503:4496] ,data[4511:4504] };
end
506 :begin
 dPIn = {data[3591:3584] ,data[3599:3592] ,data[3607:3600] ,data[3615:3608] ,data[3623:3616] ,data[3815:3808] ,data[3823:3816] ,data[3831:3824] ,data[3839:3832] ,data[3847:3840] ,data[4039:4032] ,data[4047:4040] ,data[4055:4048] ,data[4063:4056] ,data[4071:4064] ,data[4263:4256] ,data[4271:4264] ,data[4279:4272] ,data[4287:4280] ,data[4295:4288] ,data[4487:4480] ,data[4495:4488] ,data[4503:4496] ,data[4511:4504] ,data[4519:4512] };
end
507 :begin
 dPIn = {data[3599:3592] ,data[3607:3600] ,data[3615:3608] ,data[3623:3616] ,data[3631:3624] ,data[3823:3816] ,data[3831:3824] ,data[3839:3832] ,data[3847:3840] ,data[3855:3848] ,data[4047:4040] ,data[4055:4048] ,data[4063:4056] ,data[4071:4064] ,data[4079:4072] ,data[4271:4264] ,data[4279:4272] ,data[4287:4280] ,data[4295:4288] ,data[4303:4296] ,data[4495:4488] ,data[4503:4496] ,data[4511:4504] ,data[4519:4512] ,data[4527:4520] };
end
508 :begin
 dPIn = {data[3607:3600] ,data[3615:3608] ,data[3623:3616] ,data[3631:3624] ,data[3639:3632] ,data[3831:3824] ,data[3839:3832] ,data[3847:3840] ,data[3855:3848] ,data[3863:3856] ,data[4055:4048] ,data[4063:4056] ,data[4071:4064] ,data[4079:4072] ,data[4087:4080] ,data[4279:4272] ,data[4287:4280] ,data[4295:4288] ,data[4303:4296] ,data[4311:4304] ,data[4503:4496] ,data[4511:4504] ,data[4519:4512] ,data[4527:4520] ,data[4535:4528] };
end
509 :begin
 dPIn = {data[3615:3608] ,data[3623:3616] ,data[3631:3624] ,data[3639:3632] ,data[3647:3640] ,data[3839:3832] ,data[3847:3840] ,data[3855:3848] ,data[3863:3856] ,data[3871:3864] ,data[4063:4056] ,data[4071:4064] ,data[4079:4072] ,data[4087:4080] ,data[4095:4088] ,data[4287:4280] ,data[4295:4288] ,data[4303:4296] ,data[4311:4304] ,data[4319:4312] ,data[4511:4504] ,data[4519:4512] ,data[4527:4520] ,data[4535:4528] ,data[4543:4536] };
end
510 :begin
 dPIn = {data[3623:3616] ,data[3631:3624] ,data[3639:3632] ,data[3647:3640] ,data[3655:3648] ,data[3847:3840] ,data[3855:3848] ,data[3863:3856] ,data[3871:3864] ,data[3879:3872] ,data[4071:4064] ,data[4079:4072] ,data[4087:4080] ,data[4095:4088] ,data[4103:4096] ,data[4295:4288] ,data[4303:4296] ,data[4311:4304] ,data[4319:4312] ,data[4327:4320] ,data[4519:4512] ,data[4527:4520] ,data[4535:4528] ,data[4543:4536] ,data[4551:4544] };
end
511 :begin
 dPIn = {data[3631:3624] ,data[3639:3632] ,data[3647:3640] ,data[3655:3648] ,data[3663:3656] ,data[3855:3848] ,data[3863:3856] ,data[3871:3864] ,data[3879:3872] ,data[3887:3880] ,data[4079:4072] ,data[4087:4080] ,data[4095:4088] ,data[4103:4096] ,data[4111:4104] ,data[4303:4296] ,data[4311:4304] ,data[4319:4312] ,data[4327:4320] ,data[4335:4328] ,data[4527:4520] ,data[4535:4528] ,data[4543:4536] ,data[4551:4544] ,data[4559:4552] };
end
512 :begin
 dPIn = {data[3639:3632] ,data[3647:3640] ,data[3655:3648] ,data[3663:3656] ,data[3671:3664] ,data[3863:3856] ,data[3871:3864] ,data[3879:3872] ,data[3887:3880] ,data[3895:3888] ,data[4087:4080] ,data[4095:4088] ,data[4103:4096] ,data[4111:4104] ,data[4119:4112] ,data[4311:4304] ,data[4319:4312] ,data[4327:4320] ,data[4335:4328] ,data[4343:4336] ,data[4535:4528] ,data[4543:4536] ,data[4551:4544] ,data[4559:4552] ,data[4567:4560] };
end
513 :begin
 dPIn = {data[3647:3640] ,data[3655:3648] ,data[3663:3656] ,data[3671:3664] ,data[3679:3672] ,data[3871:3864] ,data[3879:3872] ,data[3887:3880] ,data[3895:3888] ,data[3903:3896] ,data[4095:4088] ,data[4103:4096] ,data[4111:4104] ,data[4119:4112] ,data[4127:4120] ,data[4319:4312] ,data[4327:4320] ,data[4335:4328] ,data[4343:4336] ,data[4351:4344] ,data[4543:4536] ,data[4551:4544] ,data[4559:4552] ,data[4567:4560] ,data[4575:4568] };
end
514 :begin
 dPIn = {data[3655:3648] ,data[3663:3656] ,data[3671:3664] ,data[3679:3672] ,data[3687:3680] ,data[3879:3872] ,data[3887:3880] ,data[3895:3888] ,data[3903:3896] ,data[3911:3904] ,data[4103:4096] ,data[4111:4104] ,data[4119:4112] ,data[4127:4120] ,data[4135:4128] ,data[4327:4320] ,data[4335:4328] ,data[4343:4336] ,data[4351:4344] ,data[4359:4352] ,data[4551:4544] ,data[4559:4552] ,data[4567:4560] ,data[4575:4568] ,data[4583:4576] };
end
515 :begin
 dPIn = {data[3663:3656] ,data[3671:3664] ,data[3679:3672] ,data[3687:3680] ,data[3695:3688] ,data[3887:3880] ,data[3895:3888] ,data[3903:3896] ,data[3911:3904] ,data[3919:3912] ,data[4111:4104] ,data[4119:4112] ,data[4127:4120] ,data[4135:4128] ,data[4143:4136] ,data[4335:4328] ,data[4343:4336] ,data[4351:4344] ,data[4359:4352] ,data[4367:4360] ,data[4559:4552] ,data[4567:4560] ,data[4575:4568] ,data[4583:4576] ,data[4591:4584] };
end
516 :begin
 dPIn = {data[3671:3664] ,data[3679:3672] ,data[3687:3680] ,data[3695:3688] ,data[3703:3696] ,data[3895:3888] ,data[3903:3896] ,data[3911:3904] ,data[3919:3912] ,data[3927:3920] ,data[4119:4112] ,data[4127:4120] ,data[4135:4128] ,data[4143:4136] ,data[4151:4144] ,data[4343:4336] ,data[4351:4344] ,data[4359:4352] ,data[4367:4360] ,data[4375:4368] ,data[4567:4560] ,data[4575:4568] ,data[4583:4576] ,data[4591:4584] ,data[4599:4592] };
end
517 :begin
 dPIn = {data[3679:3672] ,data[3687:3680] ,data[3695:3688] ,data[3703:3696] ,data[3711:3704] ,data[3903:3896] ,data[3911:3904] ,data[3919:3912] ,data[3927:3920] ,data[3935:3928] ,data[4127:4120] ,data[4135:4128] ,data[4143:4136] ,data[4151:4144] ,data[4159:4152] ,data[4351:4344] ,data[4359:4352] ,data[4367:4360] ,data[4375:4368] ,data[4383:4376] ,data[4575:4568] ,data[4583:4576] ,data[4591:4584] ,data[4599:4592] ,data[4607:4600] };
end
518 :begin
 dPIn = {data[3687:3680] ,data[3695:3688] ,data[3703:3696] ,data[3711:3704] ,data[3719:3712] ,data[3911:3904] ,data[3919:3912] ,data[3927:3920] ,data[3935:3928] ,data[3943:3936] ,data[4135:4128] ,data[4143:4136] ,data[4151:4144] ,data[4159:4152] ,data[4167:4160] ,data[4359:4352] ,data[4367:4360] ,data[4375:4368] ,data[4383:4376] ,data[4391:4384] ,data[4583:4576] ,data[4591:4584] ,data[4599:4592] ,data[4607:4600] ,data[4615:4608] };
end
519 :begin
 dPIn = {data[3695:3688] ,data[3703:3696] ,data[3711:3704] ,data[3719:3712] ,data[3727:3720] ,data[3919:3912] ,data[3927:3920] ,data[3935:3928] ,data[3943:3936] ,data[3951:3944] ,data[4143:4136] ,data[4151:4144] ,data[4159:4152] ,data[4167:4160] ,data[4175:4168] ,data[4367:4360] ,data[4375:4368] ,data[4383:4376] ,data[4391:4384] ,data[4399:4392] ,data[4591:4584] ,data[4599:4592] ,data[4607:4600] ,data[4615:4608] ,data[4623:4616] };
end
520 :begin
 dPIn = {data[3703:3696] ,data[3711:3704] ,data[3719:3712] ,data[3727:3720] ,data[3735:3728] ,data[3927:3920] ,data[3935:3928] ,data[3943:3936] ,data[3951:3944] ,data[3959:3952] ,data[4151:4144] ,data[4159:4152] ,data[4167:4160] ,data[4175:4168] ,data[4183:4176] ,data[4375:4368] ,data[4383:4376] ,data[4391:4384] ,data[4399:4392] ,data[4407:4400] ,data[4599:4592] ,data[4607:4600] ,data[4615:4608] ,data[4623:4616] ,data[4631:4624] };
end
521 :begin
 dPIn = {data[3711:3704] ,data[3719:3712] ,data[3727:3720] ,data[3735:3728] ,data[3743:3736] ,data[3935:3928] ,data[3943:3936] ,data[3951:3944] ,data[3959:3952] ,data[3967:3960] ,data[4159:4152] ,data[4167:4160] ,data[4175:4168] ,data[4183:4176] ,data[4191:4184] ,data[4383:4376] ,data[4391:4384] ,data[4399:4392] ,data[4407:4400] ,data[4415:4408] ,data[4607:4600] ,data[4615:4608] ,data[4623:4616] ,data[4631:4624] ,data[4639:4632] };
end
522 :begin
 dPIn = {data[3719:3712] ,data[3727:3720] ,data[3735:3728] ,data[3743:3736] ,data[3751:3744] ,data[3943:3936] ,data[3951:3944] ,data[3959:3952] ,data[3967:3960] ,data[3975:3968] ,data[4167:4160] ,data[4175:4168] ,data[4183:4176] ,data[4191:4184] ,data[4199:4192] ,data[4391:4384] ,data[4399:4392] ,data[4407:4400] ,data[4415:4408] ,data[4423:4416] ,data[4615:4608] ,data[4623:4616] ,data[4631:4624] ,data[4639:4632] ,data[4647:4640] };
end
523 :begin
 dPIn = {data[3727:3720] ,data[3735:3728] ,data[3743:3736] ,data[3751:3744] ,data[3759:3752] ,data[3951:3944] ,data[3959:3952] ,data[3967:3960] ,data[3975:3968] ,data[3983:3976] ,data[4175:4168] ,data[4183:4176] ,data[4191:4184] ,data[4199:4192] ,data[4207:4200] ,data[4399:4392] ,data[4407:4400] ,data[4415:4408] ,data[4423:4416] ,data[4431:4424] ,data[4623:4616] ,data[4631:4624] ,data[4639:4632] ,data[4647:4640] ,data[4655:4648] };
end
524 :begin
 dPIn = {data[3735:3728] ,data[3743:3736] ,data[3751:3744] ,data[3759:3752] ,data[3767:3760] ,data[3959:3952] ,data[3967:3960] ,data[3975:3968] ,data[3983:3976] ,data[3991:3984] ,data[4183:4176] ,data[4191:4184] ,data[4199:4192] ,data[4207:4200] ,data[4215:4208] ,data[4407:4400] ,data[4415:4408] ,data[4423:4416] ,data[4431:4424] ,data[4439:4432] ,data[4631:4624] ,data[4639:4632] ,data[4647:4640] ,data[4655:4648] ,data[4663:4656] };
end
525 :begin
 dPIn = {data[3743:3736] ,data[3751:3744] ,data[3759:3752] ,data[3767:3760] ,data[3775:3768] ,data[3967:3960] ,data[3975:3968] ,data[3983:3976] ,data[3991:3984] ,data[3999:3992] ,data[4191:4184] ,data[4199:4192] ,data[4207:4200] ,data[4215:4208] ,data[4223:4216] ,data[4415:4408] ,data[4423:4416] ,data[4431:4424] ,data[4439:4432] ,data[4447:4440] ,data[4639:4632] ,data[4647:4640] ,data[4655:4648] ,data[4663:4656] ,data[4671:4664] };
end
526 :begin
 dPIn = {data[3751:3744] ,data[3759:3752] ,data[3767:3760] ,data[3775:3768] ,data[3783:3776] ,data[3975:3968] ,data[3983:3976] ,data[3991:3984] ,data[3999:3992] ,data[4007:4000] ,data[4199:4192] ,data[4207:4200] ,data[4215:4208] ,data[4223:4216] ,data[4231:4224] ,data[4423:4416] ,data[4431:4424] ,data[4439:4432] ,data[4447:4440] ,data[4455:4448] ,data[4647:4640] ,data[4655:4648] ,data[4663:4656] ,data[4671:4664] ,data[4679:4672] };
end
527 :begin
 dPIn = {data[3759:3752] ,data[3767:3760] ,data[3775:3768] ,data[3783:3776] ,data[3791:3784] ,data[3983:3976] ,data[3991:3984] ,data[3999:3992] ,data[4007:4000] ,data[4015:4008] ,data[4207:4200] ,data[4215:4208] ,data[4223:4216] ,data[4231:4224] ,data[4239:4232] ,data[4431:4424] ,data[4439:4432] ,data[4447:4440] ,data[4455:4448] ,data[4463:4456] ,data[4655:4648] ,data[4663:4656] ,data[4671:4664] ,data[4679:4672] ,data[4687:4680] };
end
528 :begin
 dPIn = {data[3767:3760] ,data[3775:3768] ,data[3783:3776] ,data[3791:3784] ,data[3799:3792] ,data[3991:3984] ,data[3999:3992] ,data[4007:4000] ,data[4015:4008] ,data[4023:4016] ,data[4215:4208] ,data[4223:4216] ,data[4231:4224] ,data[4239:4232] ,data[4247:4240] ,data[4439:4432] ,data[4447:4440] ,data[4455:4448] ,data[4463:4456] ,data[4471:4464] ,data[4663:4656] ,data[4671:4664] ,data[4679:4672] ,data[4687:4680] ,data[4695:4688] };
end
529 :begin
 dPIn = {data[3775:3768] ,data[3783:3776] ,data[3791:3784] ,data[3799:3792] ,data[3807:3800] ,data[3999:3992] ,data[4007:4000] ,data[4015:4008] ,data[4023:4016] ,data[4031:4024] ,data[4223:4216] ,data[4231:4224] ,data[4239:4232] ,data[4247:4240] ,data[4255:4248] ,data[4447:4440] ,data[4455:4448] ,data[4463:4456] ,data[4471:4464] ,data[4479:4472] ,data[4671:4664] ,data[4679:4672] ,data[4687:4680] ,data[4695:4688] ,data[4703:4696] };
end
530 :begin
 dPIn = {data[3783:3776] ,data[3791:3784] ,data[3799:3792] ,data[3807:3800] ,0 ,data[4007:4000] ,data[4015:4008] ,data[4023:4016] ,data[4031:4024] ,0 ,data[4231:4224] ,data[4239:4232] ,data[4247:4240] ,data[4255:4248] ,0 ,data[4455:4448] ,data[4463:4456] ,data[4471:4464] ,data[4479:4472] ,0 ,data[4679:4672] ,data[4687:4680] ,data[4695:4688] ,data[4703:4696] ,0 };
end
531 :begin
 dPIn = {data[3791:3784] ,data[3799:3792] ,data[3807:3800] ,0 ,0 ,data[4015:4008] ,data[4023:4016] ,data[4031:4024] ,0 ,0 ,data[4239:4232] ,data[4247:4240] ,data[4255:4248] ,0 ,0 ,data[4463:4456] ,data[4471:4464] ,data[4479:4472] ,0 ,0 ,data[4687:4680] ,data[4695:4688] ,data[4703:4696] ,0 ,0 };
end
532 :begin
 dPIn = {0 ,0 ,data[3815:3808] ,data[3823:3816] ,data[3831:3824] ,0 ,0 ,data[4039:4032] ,data[4047:4040] ,data[4055:4048] ,0 ,0 ,data[4263:4256] ,data[4271:4264] ,data[4279:4272] ,0 ,0 ,data[4487:4480] ,data[4495:4488] ,data[4503:4496] ,0 ,0 ,data[4711:4704] ,data[4719:4712] ,data[4727:4720] };
end
533 :begin
 dPIn = {0 ,data[3815:3808] ,data[3823:3816] ,data[3831:3824] ,data[3839:3832] ,0 ,data[4039:4032] ,data[4047:4040] ,data[4055:4048] ,data[4063:4056] ,0 ,data[4263:4256] ,data[4271:4264] ,data[4279:4272] ,data[4287:4280] ,0 ,data[4487:4480] ,data[4495:4488] ,data[4503:4496] ,data[4511:4504] ,0 ,data[4711:4704] ,data[4719:4712] ,data[4727:4720] ,data[4735:4728] };
end
534 :begin
 dPIn = {data[3815:3808] ,data[3823:3816] ,data[3831:3824] ,data[3839:3832] ,data[3847:3840] ,data[4039:4032] ,data[4047:4040] ,data[4055:4048] ,data[4063:4056] ,data[4071:4064] ,data[4263:4256] ,data[4271:4264] ,data[4279:4272] ,data[4287:4280] ,data[4295:4288] ,data[4487:4480] ,data[4495:4488] ,data[4503:4496] ,data[4511:4504] ,data[4519:4512] ,data[4711:4704] ,data[4719:4712] ,data[4727:4720] ,data[4735:4728] ,data[4743:4736] };
end
535 :begin
 dPIn = {data[3823:3816] ,data[3831:3824] ,data[3839:3832] ,data[3847:3840] ,data[3855:3848] ,data[4047:4040] ,data[4055:4048] ,data[4063:4056] ,data[4071:4064] ,data[4079:4072] ,data[4271:4264] ,data[4279:4272] ,data[4287:4280] ,data[4295:4288] ,data[4303:4296] ,data[4495:4488] ,data[4503:4496] ,data[4511:4504] ,data[4519:4512] ,data[4527:4520] ,data[4719:4712] ,data[4727:4720] ,data[4735:4728] ,data[4743:4736] ,data[4751:4744] };
end
536 :begin
 dPIn = {data[3831:3824] ,data[3839:3832] ,data[3847:3840] ,data[3855:3848] ,data[3863:3856] ,data[4055:4048] ,data[4063:4056] ,data[4071:4064] ,data[4079:4072] ,data[4087:4080] ,data[4279:4272] ,data[4287:4280] ,data[4295:4288] ,data[4303:4296] ,data[4311:4304] ,data[4503:4496] ,data[4511:4504] ,data[4519:4512] ,data[4527:4520] ,data[4535:4528] ,data[4727:4720] ,data[4735:4728] ,data[4743:4736] ,data[4751:4744] ,data[4759:4752] };
end
537 :begin
 dPIn = {data[3839:3832] ,data[3847:3840] ,data[3855:3848] ,data[3863:3856] ,data[3871:3864] ,data[4063:4056] ,data[4071:4064] ,data[4079:4072] ,data[4087:4080] ,data[4095:4088] ,data[4287:4280] ,data[4295:4288] ,data[4303:4296] ,data[4311:4304] ,data[4319:4312] ,data[4511:4504] ,data[4519:4512] ,data[4527:4520] ,data[4535:4528] ,data[4543:4536] ,data[4735:4728] ,data[4743:4736] ,data[4751:4744] ,data[4759:4752] ,data[4767:4760] };
end
538 :begin
 dPIn = {data[3847:3840] ,data[3855:3848] ,data[3863:3856] ,data[3871:3864] ,data[3879:3872] ,data[4071:4064] ,data[4079:4072] ,data[4087:4080] ,data[4095:4088] ,data[4103:4096] ,data[4295:4288] ,data[4303:4296] ,data[4311:4304] ,data[4319:4312] ,data[4327:4320] ,data[4519:4512] ,data[4527:4520] ,data[4535:4528] ,data[4543:4536] ,data[4551:4544] ,data[4743:4736] ,data[4751:4744] ,data[4759:4752] ,data[4767:4760] ,data[4775:4768] };
end
539 :begin
 dPIn = {data[3855:3848] ,data[3863:3856] ,data[3871:3864] ,data[3879:3872] ,data[3887:3880] ,data[4079:4072] ,data[4087:4080] ,data[4095:4088] ,data[4103:4096] ,data[4111:4104] ,data[4303:4296] ,data[4311:4304] ,data[4319:4312] ,data[4327:4320] ,data[4335:4328] ,data[4527:4520] ,data[4535:4528] ,data[4543:4536] ,data[4551:4544] ,data[4559:4552] ,data[4751:4744] ,data[4759:4752] ,data[4767:4760] ,data[4775:4768] ,data[4783:4776] };
end
540 :begin
 dPIn = {data[3863:3856] ,data[3871:3864] ,data[3879:3872] ,data[3887:3880] ,data[3895:3888] ,data[4087:4080] ,data[4095:4088] ,data[4103:4096] ,data[4111:4104] ,data[4119:4112] ,data[4311:4304] ,data[4319:4312] ,data[4327:4320] ,data[4335:4328] ,data[4343:4336] ,data[4535:4528] ,data[4543:4536] ,data[4551:4544] ,data[4559:4552] ,data[4567:4560] ,data[4759:4752] ,data[4767:4760] ,data[4775:4768] ,data[4783:4776] ,data[4791:4784] };
end
541 :begin
 dPIn = {data[3871:3864] ,data[3879:3872] ,data[3887:3880] ,data[3895:3888] ,data[3903:3896] ,data[4095:4088] ,data[4103:4096] ,data[4111:4104] ,data[4119:4112] ,data[4127:4120] ,data[4319:4312] ,data[4327:4320] ,data[4335:4328] ,data[4343:4336] ,data[4351:4344] ,data[4543:4536] ,data[4551:4544] ,data[4559:4552] ,data[4567:4560] ,data[4575:4568] ,data[4767:4760] ,data[4775:4768] ,data[4783:4776] ,data[4791:4784] ,data[4799:4792] };
end
542 :begin
 dPIn = {data[3879:3872] ,data[3887:3880] ,data[3895:3888] ,data[3903:3896] ,data[3911:3904] ,data[4103:4096] ,data[4111:4104] ,data[4119:4112] ,data[4127:4120] ,data[4135:4128] ,data[4327:4320] ,data[4335:4328] ,data[4343:4336] ,data[4351:4344] ,data[4359:4352] ,data[4551:4544] ,data[4559:4552] ,data[4567:4560] ,data[4575:4568] ,data[4583:4576] ,data[4775:4768] ,data[4783:4776] ,data[4791:4784] ,data[4799:4792] ,data[4807:4800] };
end
543 :begin
 dPIn = {data[3887:3880] ,data[3895:3888] ,data[3903:3896] ,data[3911:3904] ,data[3919:3912] ,data[4111:4104] ,data[4119:4112] ,data[4127:4120] ,data[4135:4128] ,data[4143:4136] ,data[4335:4328] ,data[4343:4336] ,data[4351:4344] ,data[4359:4352] ,data[4367:4360] ,data[4559:4552] ,data[4567:4560] ,data[4575:4568] ,data[4583:4576] ,data[4591:4584] ,data[4783:4776] ,data[4791:4784] ,data[4799:4792] ,data[4807:4800] ,data[4815:4808] };
end
544 :begin
 dPIn = {data[3895:3888] ,data[3903:3896] ,data[3911:3904] ,data[3919:3912] ,data[3927:3920] ,data[4119:4112] ,data[4127:4120] ,data[4135:4128] ,data[4143:4136] ,data[4151:4144] ,data[4343:4336] ,data[4351:4344] ,data[4359:4352] ,data[4367:4360] ,data[4375:4368] ,data[4567:4560] ,data[4575:4568] ,data[4583:4576] ,data[4591:4584] ,data[4599:4592] ,data[4791:4784] ,data[4799:4792] ,data[4807:4800] ,data[4815:4808] ,data[4823:4816] };
end
545 :begin
 dPIn = {data[3903:3896] ,data[3911:3904] ,data[3919:3912] ,data[3927:3920] ,data[3935:3928] ,data[4127:4120] ,data[4135:4128] ,data[4143:4136] ,data[4151:4144] ,data[4159:4152] ,data[4351:4344] ,data[4359:4352] ,data[4367:4360] ,data[4375:4368] ,data[4383:4376] ,data[4575:4568] ,data[4583:4576] ,data[4591:4584] ,data[4599:4592] ,data[4607:4600] ,data[4799:4792] ,data[4807:4800] ,data[4815:4808] ,data[4823:4816] ,data[4831:4824] };
end
546 :begin
 dPIn = {data[3911:3904] ,data[3919:3912] ,data[3927:3920] ,data[3935:3928] ,data[3943:3936] ,data[4135:4128] ,data[4143:4136] ,data[4151:4144] ,data[4159:4152] ,data[4167:4160] ,data[4359:4352] ,data[4367:4360] ,data[4375:4368] ,data[4383:4376] ,data[4391:4384] ,data[4583:4576] ,data[4591:4584] ,data[4599:4592] ,data[4607:4600] ,data[4615:4608] ,data[4807:4800] ,data[4815:4808] ,data[4823:4816] ,data[4831:4824] ,data[4839:4832] };
end
547 :begin
 dPIn = {data[3919:3912] ,data[3927:3920] ,data[3935:3928] ,data[3943:3936] ,data[3951:3944] ,data[4143:4136] ,data[4151:4144] ,data[4159:4152] ,data[4167:4160] ,data[4175:4168] ,data[4367:4360] ,data[4375:4368] ,data[4383:4376] ,data[4391:4384] ,data[4399:4392] ,data[4591:4584] ,data[4599:4592] ,data[4607:4600] ,data[4615:4608] ,data[4623:4616] ,data[4815:4808] ,data[4823:4816] ,data[4831:4824] ,data[4839:4832] ,data[4847:4840] };
end
548 :begin
 dPIn = {data[3927:3920] ,data[3935:3928] ,data[3943:3936] ,data[3951:3944] ,data[3959:3952] ,data[4151:4144] ,data[4159:4152] ,data[4167:4160] ,data[4175:4168] ,data[4183:4176] ,data[4375:4368] ,data[4383:4376] ,data[4391:4384] ,data[4399:4392] ,data[4407:4400] ,data[4599:4592] ,data[4607:4600] ,data[4615:4608] ,data[4623:4616] ,data[4631:4624] ,data[4823:4816] ,data[4831:4824] ,data[4839:4832] ,data[4847:4840] ,data[4855:4848] };
end
549 :begin
 dPIn = {data[3935:3928] ,data[3943:3936] ,data[3951:3944] ,data[3959:3952] ,data[3967:3960] ,data[4159:4152] ,data[4167:4160] ,data[4175:4168] ,data[4183:4176] ,data[4191:4184] ,data[4383:4376] ,data[4391:4384] ,data[4399:4392] ,data[4407:4400] ,data[4415:4408] ,data[4607:4600] ,data[4615:4608] ,data[4623:4616] ,data[4631:4624] ,data[4639:4632] ,data[4831:4824] ,data[4839:4832] ,data[4847:4840] ,data[4855:4848] ,data[4863:4856] };
end
550 :begin
 dPIn = {data[3943:3936] ,data[3951:3944] ,data[3959:3952] ,data[3967:3960] ,data[3975:3968] ,data[4167:4160] ,data[4175:4168] ,data[4183:4176] ,data[4191:4184] ,data[4199:4192] ,data[4391:4384] ,data[4399:4392] ,data[4407:4400] ,data[4415:4408] ,data[4423:4416] ,data[4615:4608] ,data[4623:4616] ,data[4631:4624] ,data[4639:4632] ,data[4647:4640] ,data[4839:4832] ,data[4847:4840] ,data[4855:4848] ,data[4863:4856] ,data[4871:4864] };
end
551 :begin
 dPIn = {data[3951:3944] ,data[3959:3952] ,data[3967:3960] ,data[3975:3968] ,data[3983:3976] ,data[4175:4168] ,data[4183:4176] ,data[4191:4184] ,data[4199:4192] ,data[4207:4200] ,data[4399:4392] ,data[4407:4400] ,data[4415:4408] ,data[4423:4416] ,data[4431:4424] ,data[4623:4616] ,data[4631:4624] ,data[4639:4632] ,data[4647:4640] ,data[4655:4648] ,data[4847:4840] ,data[4855:4848] ,data[4863:4856] ,data[4871:4864] ,data[4879:4872] };
end
552 :begin
 dPIn = {data[3959:3952] ,data[3967:3960] ,data[3975:3968] ,data[3983:3976] ,data[3991:3984] ,data[4183:4176] ,data[4191:4184] ,data[4199:4192] ,data[4207:4200] ,data[4215:4208] ,data[4407:4400] ,data[4415:4408] ,data[4423:4416] ,data[4431:4424] ,data[4439:4432] ,data[4631:4624] ,data[4639:4632] ,data[4647:4640] ,data[4655:4648] ,data[4663:4656] ,data[4855:4848] ,data[4863:4856] ,data[4871:4864] ,data[4879:4872] ,data[4887:4880] };
end
553 :begin
 dPIn = {data[3967:3960] ,data[3975:3968] ,data[3983:3976] ,data[3991:3984] ,data[3999:3992] ,data[4191:4184] ,data[4199:4192] ,data[4207:4200] ,data[4215:4208] ,data[4223:4216] ,data[4415:4408] ,data[4423:4416] ,data[4431:4424] ,data[4439:4432] ,data[4447:4440] ,data[4639:4632] ,data[4647:4640] ,data[4655:4648] ,data[4663:4656] ,data[4671:4664] ,data[4863:4856] ,data[4871:4864] ,data[4879:4872] ,data[4887:4880] ,data[4895:4888] };
end
554 :begin
 dPIn = {data[3975:3968] ,data[3983:3976] ,data[3991:3984] ,data[3999:3992] ,data[4007:4000] ,data[4199:4192] ,data[4207:4200] ,data[4215:4208] ,data[4223:4216] ,data[4231:4224] ,data[4423:4416] ,data[4431:4424] ,data[4439:4432] ,data[4447:4440] ,data[4455:4448] ,data[4647:4640] ,data[4655:4648] ,data[4663:4656] ,data[4671:4664] ,data[4679:4672] ,data[4871:4864] ,data[4879:4872] ,data[4887:4880] ,data[4895:4888] ,data[4903:4896] };
end
555 :begin
 dPIn = {data[3983:3976] ,data[3991:3984] ,data[3999:3992] ,data[4007:4000] ,data[4015:4008] ,data[4207:4200] ,data[4215:4208] ,data[4223:4216] ,data[4231:4224] ,data[4239:4232] ,data[4431:4424] ,data[4439:4432] ,data[4447:4440] ,data[4455:4448] ,data[4463:4456] ,data[4655:4648] ,data[4663:4656] ,data[4671:4664] ,data[4679:4672] ,data[4687:4680] ,data[4879:4872] ,data[4887:4880] ,data[4895:4888] ,data[4903:4896] ,data[4911:4904] };
end
556 :begin
 dPIn = {data[3991:3984] ,data[3999:3992] ,data[4007:4000] ,data[4015:4008] ,data[4023:4016] ,data[4215:4208] ,data[4223:4216] ,data[4231:4224] ,data[4239:4232] ,data[4247:4240] ,data[4439:4432] ,data[4447:4440] ,data[4455:4448] ,data[4463:4456] ,data[4471:4464] ,data[4663:4656] ,data[4671:4664] ,data[4679:4672] ,data[4687:4680] ,data[4695:4688] ,data[4887:4880] ,data[4895:4888] ,data[4903:4896] ,data[4911:4904] ,data[4919:4912] };
end
557 :begin
 dPIn = {data[3999:3992] ,data[4007:4000] ,data[4015:4008] ,data[4023:4016] ,data[4031:4024] ,data[4223:4216] ,data[4231:4224] ,data[4239:4232] ,data[4247:4240] ,data[4255:4248] ,data[4447:4440] ,data[4455:4448] ,data[4463:4456] ,data[4471:4464] ,data[4479:4472] ,data[4671:4664] ,data[4679:4672] ,data[4687:4680] ,data[4695:4688] ,data[4703:4696] ,data[4895:4888] ,data[4903:4896] ,data[4911:4904] ,data[4919:4912] ,data[4927:4920] };
end
558 :begin
 dPIn = {data[4007:4000] ,data[4015:4008] ,data[4023:4016] ,data[4031:4024] ,0 ,data[4231:4224] ,data[4239:4232] ,data[4247:4240] ,data[4255:4248] ,0 ,data[4455:4448] ,data[4463:4456] ,data[4471:4464] ,data[4479:4472] ,0 ,data[4679:4672] ,data[4687:4680] ,data[4695:4688] ,data[4703:4696] ,0 ,data[4903:4896] ,data[4911:4904] ,data[4919:4912] ,data[4927:4920] ,0 };
end
559 :begin
 dPIn = {data[4015:4008] ,data[4023:4016] ,data[4031:4024] ,0 ,0 ,data[4239:4232] ,data[4247:4240] ,data[4255:4248] ,0 ,0 ,data[4463:4456] ,data[4471:4464] ,data[4479:4472] ,0 ,0 ,data[4687:4680] ,data[4695:4688] ,data[4703:4696] ,0 ,0 ,data[4911:4904] ,data[4919:4912] ,data[4927:4920] ,0 ,0 };
end
560 :begin
 dPIn = {0 ,0 ,data[4039:4032] ,data[4047:4040] ,data[4055:4048] ,0 ,0 ,data[4263:4256] ,data[4271:4264] ,data[4279:4272] ,0 ,0 ,data[4487:4480] ,data[4495:4488] ,data[4503:4496] ,0 ,0 ,data[4711:4704] ,data[4719:4712] ,data[4727:4720] ,0 ,0 ,data[4935:4928] ,data[4943:4936] ,data[4951:4944] };
end
561 :begin
 dPIn = {0 ,data[4039:4032] ,data[4047:4040] ,data[4055:4048] ,data[4063:4056] ,0 ,data[4263:4256] ,data[4271:4264] ,data[4279:4272] ,data[4287:4280] ,0 ,data[4487:4480] ,data[4495:4488] ,data[4503:4496] ,data[4511:4504] ,0 ,data[4711:4704] ,data[4719:4712] ,data[4727:4720] ,data[4735:4728] ,0 ,data[4935:4928] ,data[4943:4936] ,data[4951:4944] ,data[4959:4952] };
end
562 :begin
 dPIn = {data[4039:4032] ,data[4047:4040] ,data[4055:4048] ,data[4063:4056] ,data[4071:4064] ,data[4263:4256] ,data[4271:4264] ,data[4279:4272] ,data[4287:4280] ,data[4295:4288] ,data[4487:4480] ,data[4495:4488] ,data[4503:4496] ,data[4511:4504] ,data[4519:4512] ,data[4711:4704] ,data[4719:4712] ,data[4727:4720] ,data[4735:4728] ,data[4743:4736] ,data[4935:4928] ,data[4943:4936] ,data[4951:4944] ,data[4959:4952] ,data[4967:4960] };
end
563 :begin
 dPIn = {data[4047:4040] ,data[4055:4048] ,data[4063:4056] ,data[4071:4064] ,data[4079:4072] ,data[4271:4264] ,data[4279:4272] ,data[4287:4280] ,data[4295:4288] ,data[4303:4296] ,data[4495:4488] ,data[4503:4496] ,data[4511:4504] ,data[4519:4512] ,data[4527:4520] ,data[4719:4712] ,data[4727:4720] ,data[4735:4728] ,data[4743:4736] ,data[4751:4744] ,data[4943:4936] ,data[4951:4944] ,data[4959:4952] ,data[4967:4960] ,data[4975:4968] };
end
564 :begin
 dPIn = {data[4055:4048] ,data[4063:4056] ,data[4071:4064] ,data[4079:4072] ,data[4087:4080] ,data[4279:4272] ,data[4287:4280] ,data[4295:4288] ,data[4303:4296] ,data[4311:4304] ,data[4503:4496] ,data[4511:4504] ,data[4519:4512] ,data[4527:4520] ,data[4535:4528] ,data[4727:4720] ,data[4735:4728] ,data[4743:4736] ,data[4751:4744] ,data[4759:4752] ,data[4951:4944] ,data[4959:4952] ,data[4967:4960] ,data[4975:4968] ,data[4983:4976] };
end
565 :begin
 dPIn = {data[4063:4056] ,data[4071:4064] ,data[4079:4072] ,data[4087:4080] ,data[4095:4088] ,data[4287:4280] ,data[4295:4288] ,data[4303:4296] ,data[4311:4304] ,data[4319:4312] ,data[4511:4504] ,data[4519:4512] ,data[4527:4520] ,data[4535:4528] ,data[4543:4536] ,data[4735:4728] ,data[4743:4736] ,data[4751:4744] ,data[4759:4752] ,data[4767:4760] ,data[4959:4952] ,data[4967:4960] ,data[4975:4968] ,data[4983:4976] ,data[4991:4984] };
end
566 :begin
 dPIn = {data[4071:4064] ,data[4079:4072] ,data[4087:4080] ,data[4095:4088] ,data[4103:4096] ,data[4295:4288] ,data[4303:4296] ,data[4311:4304] ,data[4319:4312] ,data[4327:4320] ,data[4519:4512] ,data[4527:4520] ,data[4535:4528] ,data[4543:4536] ,data[4551:4544] ,data[4743:4736] ,data[4751:4744] ,data[4759:4752] ,data[4767:4760] ,data[4775:4768] ,data[4967:4960] ,data[4975:4968] ,data[4983:4976] ,data[4991:4984] ,data[4999:4992] };
end
567 :begin
 dPIn = {data[4079:4072] ,data[4087:4080] ,data[4095:4088] ,data[4103:4096] ,data[4111:4104] ,data[4303:4296] ,data[4311:4304] ,data[4319:4312] ,data[4327:4320] ,data[4335:4328] ,data[4527:4520] ,data[4535:4528] ,data[4543:4536] ,data[4551:4544] ,data[4559:4552] ,data[4751:4744] ,data[4759:4752] ,data[4767:4760] ,data[4775:4768] ,data[4783:4776] ,data[4975:4968] ,data[4983:4976] ,data[4991:4984] ,data[4999:4992] ,data[5007:5000] };
end
568 :begin
 dPIn = {data[4087:4080] ,data[4095:4088] ,data[4103:4096] ,data[4111:4104] ,data[4119:4112] ,data[4311:4304] ,data[4319:4312] ,data[4327:4320] ,data[4335:4328] ,data[4343:4336] ,data[4535:4528] ,data[4543:4536] ,data[4551:4544] ,data[4559:4552] ,data[4567:4560] ,data[4759:4752] ,data[4767:4760] ,data[4775:4768] ,data[4783:4776] ,data[4791:4784] ,data[4983:4976] ,data[4991:4984] ,data[4999:4992] ,data[5007:5000] ,data[5015:5008] };
end
569 :begin
 dPIn = {data[4095:4088] ,data[4103:4096] ,data[4111:4104] ,data[4119:4112] ,data[4127:4120] ,data[4319:4312] ,data[4327:4320] ,data[4335:4328] ,data[4343:4336] ,data[4351:4344] ,data[4543:4536] ,data[4551:4544] ,data[4559:4552] ,data[4567:4560] ,data[4575:4568] ,data[4767:4760] ,data[4775:4768] ,data[4783:4776] ,data[4791:4784] ,data[4799:4792] ,data[4991:4984] ,data[4999:4992] ,data[5007:5000] ,data[5015:5008] ,data[5023:5016] };
end
570 :begin
 dPIn = {data[4103:4096] ,data[4111:4104] ,data[4119:4112] ,data[4127:4120] ,data[4135:4128] ,data[4327:4320] ,data[4335:4328] ,data[4343:4336] ,data[4351:4344] ,data[4359:4352] ,data[4551:4544] ,data[4559:4552] ,data[4567:4560] ,data[4575:4568] ,data[4583:4576] ,data[4775:4768] ,data[4783:4776] ,data[4791:4784] ,data[4799:4792] ,data[4807:4800] ,data[4999:4992] ,data[5007:5000] ,data[5015:5008] ,data[5023:5016] ,data[5031:5024] };
end
571 :begin
 dPIn = {data[4111:4104] ,data[4119:4112] ,data[4127:4120] ,data[4135:4128] ,data[4143:4136] ,data[4335:4328] ,data[4343:4336] ,data[4351:4344] ,data[4359:4352] ,data[4367:4360] ,data[4559:4552] ,data[4567:4560] ,data[4575:4568] ,data[4583:4576] ,data[4591:4584] ,data[4783:4776] ,data[4791:4784] ,data[4799:4792] ,data[4807:4800] ,data[4815:4808] ,data[5007:5000] ,data[5015:5008] ,data[5023:5016] ,data[5031:5024] ,data[5039:5032] };
end
572 :begin
 dPIn = {data[4119:4112] ,data[4127:4120] ,data[4135:4128] ,data[4143:4136] ,data[4151:4144] ,data[4343:4336] ,data[4351:4344] ,data[4359:4352] ,data[4367:4360] ,data[4375:4368] ,data[4567:4560] ,data[4575:4568] ,data[4583:4576] ,data[4591:4584] ,data[4599:4592] ,data[4791:4784] ,data[4799:4792] ,data[4807:4800] ,data[4815:4808] ,data[4823:4816] ,data[5015:5008] ,data[5023:5016] ,data[5031:5024] ,data[5039:5032] ,data[5047:5040] };
end
573 :begin
 dPIn = {data[4127:4120] ,data[4135:4128] ,data[4143:4136] ,data[4151:4144] ,data[4159:4152] ,data[4351:4344] ,data[4359:4352] ,data[4367:4360] ,data[4375:4368] ,data[4383:4376] ,data[4575:4568] ,data[4583:4576] ,data[4591:4584] ,data[4599:4592] ,data[4607:4600] ,data[4799:4792] ,data[4807:4800] ,data[4815:4808] ,data[4823:4816] ,data[4831:4824] ,data[5023:5016] ,data[5031:5024] ,data[5039:5032] ,data[5047:5040] ,data[5055:5048] };
end
574 :begin
 dPIn = {data[4135:4128] ,data[4143:4136] ,data[4151:4144] ,data[4159:4152] ,data[4167:4160] ,data[4359:4352] ,data[4367:4360] ,data[4375:4368] ,data[4383:4376] ,data[4391:4384] ,data[4583:4576] ,data[4591:4584] ,data[4599:4592] ,data[4607:4600] ,data[4615:4608] ,data[4807:4800] ,data[4815:4808] ,data[4823:4816] ,data[4831:4824] ,data[4839:4832] ,data[5031:5024] ,data[5039:5032] ,data[5047:5040] ,data[5055:5048] ,data[5063:5056] };
end
575 :begin
 dPIn = {data[4143:4136] ,data[4151:4144] ,data[4159:4152] ,data[4167:4160] ,data[4175:4168] ,data[4367:4360] ,data[4375:4368] ,data[4383:4376] ,data[4391:4384] ,data[4399:4392] ,data[4591:4584] ,data[4599:4592] ,data[4607:4600] ,data[4615:4608] ,data[4623:4616] ,data[4815:4808] ,data[4823:4816] ,data[4831:4824] ,data[4839:4832] ,data[4847:4840] ,data[5039:5032] ,data[5047:5040] ,data[5055:5048] ,data[5063:5056] ,data[5071:5064] };
end
576 :begin
 dPIn = {data[4151:4144] ,data[4159:4152] ,data[4167:4160] ,data[4175:4168] ,data[4183:4176] ,data[4375:4368] ,data[4383:4376] ,data[4391:4384] ,data[4399:4392] ,data[4407:4400] ,data[4599:4592] ,data[4607:4600] ,data[4615:4608] ,data[4623:4616] ,data[4631:4624] ,data[4823:4816] ,data[4831:4824] ,data[4839:4832] ,data[4847:4840] ,data[4855:4848] ,data[5047:5040] ,data[5055:5048] ,data[5063:5056] ,data[5071:5064] ,data[5079:5072] };
end
577 :begin
 dPIn = {data[4159:4152] ,data[4167:4160] ,data[4175:4168] ,data[4183:4176] ,data[4191:4184] ,data[4383:4376] ,data[4391:4384] ,data[4399:4392] ,data[4407:4400] ,data[4415:4408] ,data[4607:4600] ,data[4615:4608] ,data[4623:4616] ,data[4631:4624] ,data[4639:4632] ,data[4831:4824] ,data[4839:4832] ,data[4847:4840] ,data[4855:4848] ,data[4863:4856] ,data[5055:5048] ,data[5063:5056] ,data[5071:5064] ,data[5079:5072] ,data[5087:5080] };
end
578 :begin
 dPIn = {data[4167:4160] ,data[4175:4168] ,data[4183:4176] ,data[4191:4184] ,data[4199:4192] ,data[4391:4384] ,data[4399:4392] ,data[4407:4400] ,data[4415:4408] ,data[4423:4416] ,data[4615:4608] ,data[4623:4616] ,data[4631:4624] ,data[4639:4632] ,data[4647:4640] ,data[4839:4832] ,data[4847:4840] ,data[4855:4848] ,data[4863:4856] ,data[4871:4864] ,data[5063:5056] ,data[5071:5064] ,data[5079:5072] ,data[5087:5080] ,data[5095:5088] };
end
579 :begin
 dPIn = {data[4175:4168] ,data[4183:4176] ,data[4191:4184] ,data[4199:4192] ,data[4207:4200] ,data[4399:4392] ,data[4407:4400] ,data[4415:4408] ,data[4423:4416] ,data[4431:4424] ,data[4623:4616] ,data[4631:4624] ,data[4639:4632] ,data[4647:4640] ,data[4655:4648] ,data[4847:4840] ,data[4855:4848] ,data[4863:4856] ,data[4871:4864] ,data[4879:4872] ,data[5071:5064] ,data[5079:5072] ,data[5087:5080] ,data[5095:5088] ,data[5103:5096] };
end
580 :begin
 dPIn = {data[4183:4176] ,data[4191:4184] ,data[4199:4192] ,data[4207:4200] ,data[4215:4208] ,data[4407:4400] ,data[4415:4408] ,data[4423:4416] ,data[4431:4424] ,data[4439:4432] ,data[4631:4624] ,data[4639:4632] ,data[4647:4640] ,data[4655:4648] ,data[4663:4656] ,data[4855:4848] ,data[4863:4856] ,data[4871:4864] ,data[4879:4872] ,data[4887:4880] ,data[5079:5072] ,data[5087:5080] ,data[5095:5088] ,data[5103:5096] ,data[5111:5104] };
end
581 :begin
 dPIn = {data[4191:4184] ,data[4199:4192] ,data[4207:4200] ,data[4215:4208] ,data[4223:4216] ,data[4415:4408] ,data[4423:4416] ,data[4431:4424] ,data[4439:4432] ,data[4447:4440] ,data[4639:4632] ,data[4647:4640] ,data[4655:4648] ,data[4663:4656] ,data[4671:4664] ,data[4863:4856] ,data[4871:4864] ,data[4879:4872] ,data[4887:4880] ,data[4895:4888] ,data[5087:5080] ,data[5095:5088] ,data[5103:5096] ,data[5111:5104] ,data[5119:5112] };
end
582 :begin
 dPIn = {data[4199:4192] ,data[4207:4200] ,data[4215:4208] ,data[4223:4216] ,data[4231:4224] ,data[4423:4416] ,data[4431:4424] ,data[4439:4432] ,data[4447:4440] ,data[4455:4448] ,data[4647:4640] ,data[4655:4648] ,data[4663:4656] ,data[4671:4664] ,data[4679:4672] ,data[4871:4864] ,data[4879:4872] ,data[4887:4880] ,data[4895:4888] ,data[4903:4896] ,data[5095:5088] ,data[5103:5096] ,data[5111:5104] ,data[5119:5112] ,data[5127:5120] };
end
583 :begin
 dPIn = {data[4207:4200] ,data[4215:4208] ,data[4223:4216] ,data[4231:4224] ,data[4239:4232] ,data[4431:4424] ,data[4439:4432] ,data[4447:4440] ,data[4455:4448] ,data[4463:4456] ,data[4655:4648] ,data[4663:4656] ,data[4671:4664] ,data[4679:4672] ,data[4687:4680] ,data[4879:4872] ,data[4887:4880] ,data[4895:4888] ,data[4903:4896] ,data[4911:4904] ,data[5103:5096] ,data[5111:5104] ,data[5119:5112] ,data[5127:5120] ,data[5135:5128] };
end
584 :begin
 dPIn = {data[4215:4208] ,data[4223:4216] ,data[4231:4224] ,data[4239:4232] ,data[4247:4240] ,data[4439:4432] ,data[4447:4440] ,data[4455:4448] ,data[4463:4456] ,data[4471:4464] ,data[4663:4656] ,data[4671:4664] ,data[4679:4672] ,data[4687:4680] ,data[4695:4688] ,data[4887:4880] ,data[4895:4888] ,data[4903:4896] ,data[4911:4904] ,data[4919:4912] ,data[5111:5104] ,data[5119:5112] ,data[5127:5120] ,data[5135:5128] ,data[5143:5136] };
end
585 :begin
 dPIn = {data[4223:4216] ,data[4231:4224] ,data[4239:4232] ,data[4247:4240] ,data[4255:4248] ,data[4447:4440] ,data[4455:4448] ,data[4463:4456] ,data[4471:4464] ,data[4479:4472] ,data[4671:4664] ,data[4679:4672] ,data[4687:4680] ,data[4695:4688] ,data[4703:4696] ,data[4895:4888] ,data[4903:4896] ,data[4911:4904] ,data[4919:4912] ,data[4927:4920] ,data[5119:5112] ,data[5127:5120] ,data[5135:5128] ,data[5143:5136] ,data[5151:5144] };
end
586 :begin
 dPIn = {data[4231:4224] ,data[4239:4232] ,data[4247:4240] ,data[4255:4248] ,0 ,data[4455:4448] ,data[4463:4456] ,data[4471:4464] ,data[4479:4472] ,0 ,data[4679:4672] ,data[4687:4680] ,data[4695:4688] ,data[4703:4696] ,0 ,data[4903:4896] ,data[4911:4904] ,data[4919:4912] ,data[4927:4920] ,0 ,data[5127:5120] ,data[5135:5128] ,data[5143:5136] ,data[5151:5144] ,0 };
end
587 :begin
 dPIn = {data[4239:4232] ,data[4247:4240] ,data[4255:4248] ,0 ,0 ,data[4463:4456] ,data[4471:4464] ,data[4479:4472] ,0 ,0 ,data[4687:4680] ,data[4695:4688] ,data[4703:4696] ,0 ,0 ,data[4911:4904] ,data[4919:4912] ,data[4927:4920] ,0 ,0 ,data[5135:5128] ,data[5143:5136] ,data[5151:5144] ,0 ,0 };
end
588 :begin
 dPIn = {0 ,0 ,data[4263:4256] ,data[4271:4264] ,data[4279:4272] ,0 ,0 ,data[4487:4480] ,data[4495:4488] ,data[4503:4496] ,0 ,0 ,data[4711:4704] ,data[4719:4712] ,data[4727:4720] ,0 ,0 ,data[4935:4928] ,data[4943:4936] ,data[4951:4944] ,0 ,0 ,data[5159:5152] ,data[5167:5160] ,data[5175:5168] };
end
589 :begin
 dPIn = {0 ,data[4263:4256] ,data[4271:4264] ,data[4279:4272] ,data[4287:4280] ,0 ,data[4487:4480] ,data[4495:4488] ,data[4503:4496] ,data[4511:4504] ,0 ,data[4711:4704] ,data[4719:4712] ,data[4727:4720] ,data[4735:4728] ,0 ,data[4935:4928] ,data[4943:4936] ,data[4951:4944] ,data[4959:4952] ,0 ,data[5159:5152] ,data[5167:5160] ,data[5175:5168] ,data[5183:5176] };
end
590 :begin
 dPIn = {data[4263:4256] ,data[4271:4264] ,data[4279:4272] ,data[4287:4280] ,data[4295:4288] ,data[4487:4480] ,data[4495:4488] ,data[4503:4496] ,data[4511:4504] ,data[4519:4512] ,data[4711:4704] ,data[4719:4712] ,data[4727:4720] ,data[4735:4728] ,data[4743:4736] ,data[4935:4928] ,data[4943:4936] ,data[4951:4944] ,data[4959:4952] ,data[4967:4960] ,data[5159:5152] ,data[5167:5160] ,data[5175:5168] ,data[5183:5176] ,data[5191:5184] };
end
591 :begin
 dPIn = {data[4271:4264] ,data[4279:4272] ,data[4287:4280] ,data[4295:4288] ,data[4303:4296] ,data[4495:4488] ,data[4503:4496] ,data[4511:4504] ,data[4519:4512] ,data[4527:4520] ,data[4719:4712] ,data[4727:4720] ,data[4735:4728] ,data[4743:4736] ,data[4751:4744] ,data[4943:4936] ,data[4951:4944] ,data[4959:4952] ,data[4967:4960] ,data[4975:4968] ,data[5167:5160] ,data[5175:5168] ,data[5183:5176] ,data[5191:5184] ,data[5199:5192] };
end
592 :begin
 dPIn = {data[4279:4272] ,data[4287:4280] ,data[4295:4288] ,data[4303:4296] ,data[4311:4304] ,data[4503:4496] ,data[4511:4504] ,data[4519:4512] ,data[4527:4520] ,data[4535:4528] ,data[4727:4720] ,data[4735:4728] ,data[4743:4736] ,data[4751:4744] ,data[4759:4752] ,data[4951:4944] ,data[4959:4952] ,data[4967:4960] ,data[4975:4968] ,data[4983:4976] ,data[5175:5168] ,data[5183:5176] ,data[5191:5184] ,data[5199:5192] ,data[5207:5200] };
end
593 :begin
 dPIn = {data[4287:4280] ,data[4295:4288] ,data[4303:4296] ,data[4311:4304] ,data[4319:4312] ,data[4511:4504] ,data[4519:4512] ,data[4527:4520] ,data[4535:4528] ,data[4543:4536] ,data[4735:4728] ,data[4743:4736] ,data[4751:4744] ,data[4759:4752] ,data[4767:4760] ,data[4959:4952] ,data[4967:4960] ,data[4975:4968] ,data[4983:4976] ,data[4991:4984] ,data[5183:5176] ,data[5191:5184] ,data[5199:5192] ,data[5207:5200] ,data[5215:5208] };
end
594 :begin
 dPIn = {data[4295:4288] ,data[4303:4296] ,data[4311:4304] ,data[4319:4312] ,data[4327:4320] ,data[4519:4512] ,data[4527:4520] ,data[4535:4528] ,data[4543:4536] ,data[4551:4544] ,data[4743:4736] ,data[4751:4744] ,data[4759:4752] ,data[4767:4760] ,data[4775:4768] ,data[4967:4960] ,data[4975:4968] ,data[4983:4976] ,data[4991:4984] ,data[4999:4992] ,data[5191:5184] ,data[5199:5192] ,data[5207:5200] ,data[5215:5208] ,data[5223:5216] };
end
595 :begin
 dPIn = {data[4303:4296] ,data[4311:4304] ,data[4319:4312] ,data[4327:4320] ,data[4335:4328] ,data[4527:4520] ,data[4535:4528] ,data[4543:4536] ,data[4551:4544] ,data[4559:4552] ,data[4751:4744] ,data[4759:4752] ,data[4767:4760] ,data[4775:4768] ,data[4783:4776] ,data[4975:4968] ,data[4983:4976] ,data[4991:4984] ,data[4999:4992] ,data[5007:5000] ,data[5199:5192] ,data[5207:5200] ,data[5215:5208] ,data[5223:5216] ,data[5231:5224] };
end
596 :begin
 dPIn = {data[4311:4304] ,data[4319:4312] ,data[4327:4320] ,data[4335:4328] ,data[4343:4336] ,data[4535:4528] ,data[4543:4536] ,data[4551:4544] ,data[4559:4552] ,data[4567:4560] ,data[4759:4752] ,data[4767:4760] ,data[4775:4768] ,data[4783:4776] ,data[4791:4784] ,data[4983:4976] ,data[4991:4984] ,data[4999:4992] ,data[5007:5000] ,data[5015:5008] ,data[5207:5200] ,data[5215:5208] ,data[5223:5216] ,data[5231:5224] ,data[5239:5232] };
end
597 :begin
 dPIn = {data[4319:4312] ,data[4327:4320] ,data[4335:4328] ,data[4343:4336] ,data[4351:4344] ,data[4543:4536] ,data[4551:4544] ,data[4559:4552] ,data[4567:4560] ,data[4575:4568] ,data[4767:4760] ,data[4775:4768] ,data[4783:4776] ,data[4791:4784] ,data[4799:4792] ,data[4991:4984] ,data[4999:4992] ,data[5007:5000] ,data[5015:5008] ,data[5023:5016] ,data[5215:5208] ,data[5223:5216] ,data[5231:5224] ,data[5239:5232] ,data[5247:5240] };
end
598 :begin
 dPIn = {data[4327:4320] ,data[4335:4328] ,data[4343:4336] ,data[4351:4344] ,data[4359:4352] ,data[4551:4544] ,data[4559:4552] ,data[4567:4560] ,data[4575:4568] ,data[4583:4576] ,data[4775:4768] ,data[4783:4776] ,data[4791:4784] ,data[4799:4792] ,data[4807:4800] ,data[4999:4992] ,data[5007:5000] ,data[5015:5008] ,data[5023:5016] ,data[5031:5024] ,data[5223:5216] ,data[5231:5224] ,data[5239:5232] ,data[5247:5240] ,data[5255:5248] };
end
599 :begin
 dPIn = {data[4335:4328] ,data[4343:4336] ,data[4351:4344] ,data[4359:4352] ,data[4367:4360] ,data[4559:4552] ,data[4567:4560] ,data[4575:4568] ,data[4583:4576] ,data[4591:4584] ,data[4783:4776] ,data[4791:4784] ,data[4799:4792] ,data[4807:4800] ,data[4815:4808] ,data[5007:5000] ,data[5015:5008] ,data[5023:5016] ,data[5031:5024] ,data[5039:5032] ,data[5231:5224] ,data[5239:5232] ,data[5247:5240] ,data[5255:5248] ,data[5263:5256] };
end
600 :begin
 dPIn = {data[4343:4336] ,data[4351:4344] ,data[4359:4352] ,data[4367:4360] ,data[4375:4368] ,data[4567:4560] ,data[4575:4568] ,data[4583:4576] ,data[4591:4584] ,data[4599:4592] ,data[4791:4784] ,data[4799:4792] ,data[4807:4800] ,data[4815:4808] ,data[4823:4816] ,data[5015:5008] ,data[5023:5016] ,data[5031:5024] ,data[5039:5032] ,data[5047:5040] ,data[5239:5232] ,data[5247:5240] ,data[5255:5248] ,data[5263:5256] ,data[5271:5264] };
end
601 :begin
 dPIn = {data[4351:4344] ,data[4359:4352] ,data[4367:4360] ,data[4375:4368] ,data[4383:4376] ,data[4575:4568] ,data[4583:4576] ,data[4591:4584] ,data[4599:4592] ,data[4607:4600] ,data[4799:4792] ,data[4807:4800] ,data[4815:4808] ,data[4823:4816] ,data[4831:4824] ,data[5023:5016] ,data[5031:5024] ,data[5039:5032] ,data[5047:5040] ,data[5055:5048] ,data[5247:5240] ,data[5255:5248] ,data[5263:5256] ,data[5271:5264] ,data[5279:5272] };
end
602 :begin
 dPIn = {data[4359:4352] ,data[4367:4360] ,data[4375:4368] ,data[4383:4376] ,data[4391:4384] ,data[4583:4576] ,data[4591:4584] ,data[4599:4592] ,data[4607:4600] ,data[4615:4608] ,data[4807:4800] ,data[4815:4808] ,data[4823:4816] ,data[4831:4824] ,data[4839:4832] ,data[5031:5024] ,data[5039:5032] ,data[5047:5040] ,data[5055:5048] ,data[5063:5056] ,data[5255:5248] ,data[5263:5256] ,data[5271:5264] ,data[5279:5272] ,data[5287:5280] };
end
603 :begin
 dPIn = {data[4367:4360] ,data[4375:4368] ,data[4383:4376] ,data[4391:4384] ,data[4399:4392] ,data[4591:4584] ,data[4599:4592] ,data[4607:4600] ,data[4615:4608] ,data[4623:4616] ,data[4815:4808] ,data[4823:4816] ,data[4831:4824] ,data[4839:4832] ,data[4847:4840] ,data[5039:5032] ,data[5047:5040] ,data[5055:5048] ,data[5063:5056] ,data[5071:5064] ,data[5263:5256] ,data[5271:5264] ,data[5279:5272] ,data[5287:5280] ,data[5295:5288] };
end
604 :begin
 dPIn = {data[4375:4368] ,data[4383:4376] ,data[4391:4384] ,data[4399:4392] ,data[4407:4400] ,data[4599:4592] ,data[4607:4600] ,data[4615:4608] ,data[4623:4616] ,data[4631:4624] ,data[4823:4816] ,data[4831:4824] ,data[4839:4832] ,data[4847:4840] ,data[4855:4848] ,data[5047:5040] ,data[5055:5048] ,data[5063:5056] ,data[5071:5064] ,data[5079:5072] ,data[5271:5264] ,data[5279:5272] ,data[5287:5280] ,data[5295:5288] ,data[5303:5296] };
end
605 :begin
 dPIn = {data[4383:4376] ,data[4391:4384] ,data[4399:4392] ,data[4407:4400] ,data[4415:4408] ,data[4607:4600] ,data[4615:4608] ,data[4623:4616] ,data[4631:4624] ,data[4639:4632] ,data[4831:4824] ,data[4839:4832] ,data[4847:4840] ,data[4855:4848] ,data[4863:4856] ,data[5055:5048] ,data[5063:5056] ,data[5071:5064] ,data[5079:5072] ,data[5087:5080] ,data[5279:5272] ,data[5287:5280] ,data[5295:5288] ,data[5303:5296] ,data[5311:5304] };
end
606 :begin
 dPIn = {data[4391:4384] ,data[4399:4392] ,data[4407:4400] ,data[4415:4408] ,data[4423:4416] ,data[4615:4608] ,data[4623:4616] ,data[4631:4624] ,data[4639:4632] ,data[4647:4640] ,data[4839:4832] ,data[4847:4840] ,data[4855:4848] ,data[4863:4856] ,data[4871:4864] ,data[5063:5056] ,data[5071:5064] ,data[5079:5072] ,data[5087:5080] ,data[5095:5088] ,data[5287:5280] ,data[5295:5288] ,data[5303:5296] ,data[5311:5304] ,data[5319:5312] };
end
607 :begin
 dPIn = {data[4399:4392] ,data[4407:4400] ,data[4415:4408] ,data[4423:4416] ,data[4431:4424] ,data[4623:4616] ,data[4631:4624] ,data[4639:4632] ,data[4647:4640] ,data[4655:4648] ,data[4847:4840] ,data[4855:4848] ,data[4863:4856] ,data[4871:4864] ,data[4879:4872] ,data[5071:5064] ,data[5079:5072] ,data[5087:5080] ,data[5095:5088] ,data[5103:5096] ,data[5295:5288] ,data[5303:5296] ,data[5311:5304] ,data[5319:5312] ,data[5327:5320] };
end
608 :begin
 dPIn = {data[4407:4400] ,data[4415:4408] ,data[4423:4416] ,data[4431:4424] ,data[4439:4432] ,data[4631:4624] ,data[4639:4632] ,data[4647:4640] ,data[4655:4648] ,data[4663:4656] ,data[4855:4848] ,data[4863:4856] ,data[4871:4864] ,data[4879:4872] ,data[4887:4880] ,data[5079:5072] ,data[5087:5080] ,data[5095:5088] ,data[5103:5096] ,data[5111:5104] ,data[5303:5296] ,data[5311:5304] ,data[5319:5312] ,data[5327:5320] ,data[5335:5328] };
end
609 :begin
 dPIn = {data[4415:4408] ,data[4423:4416] ,data[4431:4424] ,data[4439:4432] ,data[4447:4440] ,data[4639:4632] ,data[4647:4640] ,data[4655:4648] ,data[4663:4656] ,data[4671:4664] ,data[4863:4856] ,data[4871:4864] ,data[4879:4872] ,data[4887:4880] ,data[4895:4888] ,data[5087:5080] ,data[5095:5088] ,data[5103:5096] ,data[5111:5104] ,data[5119:5112] ,data[5311:5304] ,data[5319:5312] ,data[5327:5320] ,data[5335:5328] ,data[5343:5336] };
end
610 :begin
 dPIn = {data[4423:4416] ,data[4431:4424] ,data[4439:4432] ,data[4447:4440] ,data[4455:4448] ,data[4647:4640] ,data[4655:4648] ,data[4663:4656] ,data[4671:4664] ,data[4679:4672] ,data[4871:4864] ,data[4879:4872] ,data[4887:4880] ,data[4895:4888] ,data[4903:4896] ,data[5095:5088] ,data[5103:5096] ,data[5111:5104] ,data[5119:5112] ,data[5127:5120] ,data[5319:5312] ,data[5327:5320] ,data[5335:5328] ,data[5343:5336] ,data[5351:5344] };
end
611 :begin
 dPIn = {data[4431:4424] ,data[4439:4432] ,data[4447:4440] ,data[4455:4448] ,data[4463:4456] ,data[4655:4648] ,data[4663:4656] ,data[4671:4664] ,data[4679:4672] ,data[4687:4680] ,data[4879:4872] ,data[4887:4880] ,data[4895:4888] ,data[4903:4896] ,data[4911:4904] ,data[5103:5096] ,data[5111:5104] ,data[5119:5112] ,data[5127:5120] ,data[5135:5128] ,data[5327:5320] ,data[5335:5328] ,data[5343:5336] ,data[5351:5344] ,data[5359:5352] };
end
612 :begin
 dPIn = {data[4439:4432] ,data[4447:4440] ,data[4455:4448] ,data[4463:4456] ,data[4471:4464] ,data[4663:4656] ,data[4671:4664] ,data[4679:4672] ,data[4687:4680] ,data[4695:4688] ,data[4887:4880] ,data[4895:4888] ,data[4903:4896] ,data[4911:4904] ,data[4919:4912] ,data[5111:5104] ,data[5119:5112] ,data[5127:5120] ,data[5135:5128] ,data[5143:5136] ,data[5335:5328] ,data[5343:5336] ,data[5351:5344] ,data[5359:5352] ,data[5367:5360] };
end
613 :begin
 dPIn = {data[4447:4440] ,data[4455:4448] ,data[4463:4456] ,data[4471:4464] ,data[4479:4472] ,data[4671:4664] ,data[4679:4672] ,data[4687:4680] ,data[4695:4688] ,data[4703:4696] ,data[4895:4888] ,data[4903:4896] ,data[4911:4904] ,data[4919:4912] ,data[4927:4920] ,data[5119:5112] ,data[5127:5120] ,data[5135:5128] ,data[5143:5136] ,data[5151:5144] ,data[5343:5336] ,data[5351:5344] ,data[5359:5352] ,data[5367:5360] ,data[5375:5368] };
end
614 :begin
 dPIn = {data[4455:4448] ,data[4463:4456] ,data[4471:4464] ,data[4479:4472] ,0 ,data[4679:4672] ,data[4687:4680] ,data[4695:4688] ,data[4703:4696] ,0 ,data[4903:4896] ,data[4911:4904] ,data[4919:4912] ,data[4927:4920] ,0 ,data[5127:5120] ,data[5135:5128] ,data[5143:5136] ,data[5151:5144] ,0 ,data[5351:5344] ,data[5359:5352] ,data[5367:5360] ,data[5375:5368] ,0 };
end
615 :begin
 dPIn = {data[4463:4456] ,data[4471:4464] ,data[4479:4472] ,0 ,0 ,data[4687:4680] ,data[4695:4688] ,data[4703:4696] ,0 ,0 ,data[4911:4904] ,data[4919:4912] ,data[4927:4920] ,0 ,0 ,data[5135:5128] ,data[5143:5136] ,data[5151:5144] ,0 ,0 ,data[5359:5352] ,data[5367:5360] ,data[5375:5368] ,0 ,0 };
end
616 :begin
 dPIn = {0 ,0 ,data[4487:4480] ,data[4495:4488] ,data[4503:4496] ,0 ,0 ,data[4711:4704] ,data[4719:4712] ,data[4727:4720] ,0 ,0 ,data[4935:4928] ,data[4943:4936] ,data[4951:4944] ,0 ,0 ,data[5159:5152] ,data[5167:5160] ,data[5175:5168] ,0 ,0 ,data[5383:5376] ,data[5391:5384] ,data[5399:5392] };
end
617 :begin
 dPIn = {0 ,data[4487:4480] ,data[4495:4488] ,data[4503:4496] ,data[4511:4504] ,0 ,data[4711:4704] ,data[4719:4712] ,data[4727:4720] ,data[4735:4728] ,0 ,data[4935:4928] ,data[4943:4936] ,data[4951:4944] ,data[4959:4952] ,0 ,data[5159:5152] ,data[5167:5160] ,data[5175:5168] ,data[5183:5176] ,0 ,data[5383:5376] ,data[5391:5384] ,data[5399:5392] ,data[5407:5400] };
end
618 :begin
 dPIn = {data[4487:4480] ,data[4495:4488] ,data[4503:4496] ,data[4511:4504] ,data[4519:4512] ,data[4711:4704] ,data[4719:4712] ,data[4727:4720] ,data[4735:4728] ,data[4743:4736] ,data[4935:4928] ,data[4943:4936] ,data[4951:4944] ,data[4959:4952] ,data[4967:4960] ,data[5159:5152] ,data[5167:5160] ,data[5175:5168] ,data[5183:5176] ,data[5191:5184] ,data[5383:5376] ,data[5391:5384] ,data[5399:5392] ,data[5407:5400] ,data[5415:5408] };
end
619 :begin
 dPIn = {data[4495:4488] ,data[4503:4496] ,data[4511:4504] ,data[4519:4512] ,data[4527:4520] ,data[4719:4712] ,data[4727:4720] ,data[4735:4728] ,data[4743:4736] ,data[4751:4744] ,data[4943:4936] ,data[4951:4944] ,data[4959:4952] ,data[4967:4960] ,data[4975:4968] ,data[5167:5160] ,data[5175:5168] ,data[5183:5176] ,data[5191:5184] ,data[5199:5192] ,data[5391:5384] ,data[5399:5392] ,data[5407:5400] ,data[5415:5408] ,data[5423:5416] };
end
620 :begin
 dPIn = {data[4503:4496] ,data[4511:4504] ,data[4519:4512] ,data[4527:4520] ,data[4535:4528] ,data[4727:4720] ,data[4735:4728] ,data[4743:4736] ,data[4751:4744] ,data[4759:4752] ,data[4951:4944] ,data[4959:4952] ,data[4967:4960] ,data[4975:4968] ,data[4983:4976] ,data[5175:5168] ,data[5183:5176] ,data[5191:5184] ,data[5199:5192] ,data[5207:5200] ,data[5399:5392] ,data[5407:5400] ,data[5415:5408] ,data[5423:5416] ,data[5431:5424] };
end
621 :begin
 dPIn = {data[4511:4504] ,data[4519:4512] ,data[4527:4520] ,data[4535:4528] ,data[4543:4536] ,data[4735:4728] ,data[4743:4736] ,data[4751:4744] ,data[4759:4752] ,data[4767:4760] ,data[4959:4952] ,data[4967:4960] ,data[4975:4968] ,data[4983:4976] ,data[4991:4984] ,data[5183:5176] ,data[5191:5184] ,data[5199:5192] ,data[5207:5200] ,data[5215:5208] ,data[5407:5400] ,data[5415:5408] ,data[5423:5416] ,data[5431:5424] ,data[5439:5432] };
end
622 :begin
 dPIn = {data[4519:4512] ,data[4527:4520] ,data[4535:4528] ,data[4543:4536] ,data[4551:4544] ,data[4743:4736] ,data[4751:4744] ,data[4759:4752] ,data[4767:4760] ,data[4775:4768] ,data[4967:4960] ,data[4975:4968] ,data[4983:4976] ,data[4991:4984] ,data[4999:4992] ,data[5191:5184] ,data[5199:5192] ,data[5207:5200] ,data[5215:5208] ,data[5223:5216] ,data[5415:5408] ,data[5423:5416] ,data[5431:5424] ,data[5439:5432] ,data[5447:5440] };
end
623 :begin
 dPIn = {data[4527:4520] ,data[4535:4528] ,data[4543:4536] ,data[4551:4544] ,data[4559:4552] ,data[4751:4744] ,data[4759:4752] ,data[4767:4760] ,data[4775:4768] ,data[4783:4776] ,data[4975:4968] ,data[4983:4976] ,data[4991:4984] ,data[4999:4992] ,data[5007:5000] ,data[5199:5192] ,data[5207:5200] ,data[5215:5208] ,data[5223:5216] ,data[5231:5224] ,data[5423:5416] ,data[5431:5424] ,data[5439:5432] ,data[5447:5440] ,data[5455:5448] };
end
624 :begin
 dPIn = {data[4535:4528] ,data[4543:4536] ,data[4551:4544] ,data[4559:4552] ,data[4567:4560] ,data[4759:4752] ,data[4767:4760] ,data[4775:4768] ,data[4783:4776] ,data[4791:4784] ,data[4983:4976] ,data[4991:4984] ,data[4999:4992] ,data[5007:5000] ,data[5015:5008] ,data[5207:5200] ,data[5215:5208] ,data[5223:5216] ,data[5231:5224] ,data[5239:5232] ,data[5431:5424] ,data[5439:5432] ,data[5447:5440] ,data[5455:5448] ,data[5463:5456] };
end
625 :begin
 dPIn = {data[4543:4536] ,data[4551:4544] ,data[4559:4552] ,data[4567:4560] ,data[4575:4568] ,data[4767:4760] ,data[4775:4768] ,data[4783:4776] ,data[4791:4784] ,data[4799:4792] ,data[4991:4984] ,data[4999:4992] ,data[5007:5000] ,data[5015:5008] ,data[5023:5016] ,data[5215:5208] ,data[5223:5216] ,data[5231:5224] ,data[5239:5232] ,data[5247:5240] ,data[5439:5432] ,data[5447:5440] ,data[5455:5448] ,data[5463:5456] ,data[5471:5464] };
end
626 :begin
 dPIn = {data[4551:4544] ,data[4559:4552] ,data[4567:4560] ,data[4575:4568] ,data[4583:4576] ,data[4775:4768] ,data[4783:4776] ,data[4791:4784] ,data[4799:4792] ,data[4807:4800] ,data[4999:4992] ,data[5007:5000] ,data[5015:5008] ,data[5023:5016] ,data[5031:5024] ,data[5223:5216] ,data[5231:5224] ,data[5239:5232] ,data[5247:5240] ,data[5255:5248] ,data[5447:5440] ,data[5455:5448] ,data[5463:5456] ,data[5471:5464] ,data[5479:5472] };
end
627 :begin
 dPIn = {data[4559:4552] ,data[4567:4560] ,data[4575:4568] ,data[4583:4576] ,data[4591:4584] ,data[4783:4776] ,data[4791:4784] ,data[4799:4792] ,data[4807:4800] ,data[4815:4808] ,data[5007:5000] ,data[5015:5008] ,data[5023:5016] ,data[5031:5024] ,data[5039:5032] ,data[5231:5224] ,data[5239:5232] ,data[5247:5240] ,data[5255:5248] ,data[5263:5256] ,data[5455:5448] ,data[5463:5456] ,data[5471:5464] ,data[5479:5472] ,data[5487:5480] };
end
628 :begin
 dPIn = {data[4567:4560] ,data[4575:4568] ,data[4583:4576] ,data[4591:4584] ,data[4599:4592] ,data[4791:4784] ,data[4799:4792] ,data[4807:4800] ,data[4815:4808] ,data[4823:4816] ,data[5015:5008] ,data[5023:5016] ,data[5031:5024] ,data[5039:5032] ,data[5047:5040] ,data[5239:5232] ,data[5247:5240] ,data[5255:5248] ,data[5263:5256] ,data[5271:5264] ,data[5463:5456] ,data[5471:5464] ,data[5479:5472] ,data[5487:5480] ,data[5495:5488] };
end
629 :begin
 dPIn = {data[4575:4568] ,data[4583:4576] ,data[4591:4584] ,data[4599:4592] ,data[4607:4600] ,data[4799:4792] ,data[4807:4800] ,data[4815:4808] ,data[4823:4816] ,data[4831:4824] ,data[5023:5016] ,data[5031:5024] ,data[5039:5032] ,data[5047:5040] ,data[5055:5048] ,data[5247:5240] ,data[5255:5248] ,data[5263:5256] ,data[5271:5264] ,data[5279:5272] ,data[5471:5464] ,data[5479:5472] ,data[5487:5480] ,data[5495:5488] ,data[5503:5496] };
end
630 :begin
 dPIn = {data[4583:4576] ,data[4591:4584] ,data[4599:4592] ,data[4607:4600] ,data[4615:4608] ,data[4807:4800] ,data[4815:4808] ,data[4823:4816] ,data[4831:4824] ,data[4839:4832] ,data[5031:5024] ,data[5039:5032] ,data[5047:5040] ,data[5055:5048] ,data[5063:5056] ,data[5255:5248] ,data[5263:5256] ,data[5271:5264] ,data[5279:5272] ,data[5287:5280] ,data[5479:5472] ,data[5487:5480] ,data[5495:5488] ,data[5503:5496] ,data[5511:5504] };
end
631 :begin
 dPIn = {data[4591:4584] ,data[4599:4592] ,data[4607:4600] ,data[4615:4608] ,data[4623:4616] ,data[4815:4808] ,data[4823:4816] ,data[4831:4824] ,data[4839:4832] ,data[4847:4840] ,data[5039:5032] ,data[5047:5040] ,data[5055:5048] ,data[5063:5056] ,data[5071:5064] ,data[5263:5256] ,data[5271:5264] ,data[5279:5272] ,data[5287:5280] ,data[5295:5288] ,data[5487:5480] ,data[5495:5488] ,data[5503:5496] ,data[5511:5504] ,data[5519:5512] };
end
632 :begin
 dPIn = {data[4599:4592] ,data[4607:4600] ,data[4615:4608] ,data[4623:4616] ,data[4631:4624] ,data[4823:4816] ,data[4831:4824] ,data[4839:4832] ,data[4847:4840] ,data[4855:4848] ,data[5047:5040] ,data[5055:5048] ,data[5063:5056] ,data[5071:5064] ,data[5079:5072] ,data[5271:5264] ,data[5279:5272] ,data[5287:5280] ,data[5295:5288] ,data[5303:5296] ,data[5495:5488] ,data[5503:5496] ,data[5511:5504] ,data[5519:5512] ,data[5527:5520] };
end
633 :begin
 dPIn = {data[4607:4600] ,data[4615:4608] ,data[4623:4616] ,data[4631:4624] ,data[4639:4632] ,data[4831:4824] ,data[4839:4832] ,data[4847:4840] ,data[4855:4848] ,data[4863:4856] ,data[5055:5048] ,data[5063:5056] ,data[5071:5064] ,data[5079:5072] ,data[5087:5080] ,data[5279:5272] ,data[5287:5280] ,data[5295:5288] ,data[5303:5296] ,data[5311:5304] ,data[5503:5496] ,data[5511:5504] ,data[5519:5512] ,data[5527:5520] ,data[5535:5528] };
end
634 :begin
 dPIn = {data[4615:4608] ,data[4623:4616] ,data[4631:4624] ,data[4639:4632] ,data[4647:4640] ,data[4839:4832] ,data[4847:4840] ,data[4855:4848] ,data[4863:4856] ,data[4871:4864] ,data[5063:5056] ,data[5071:5064] ,data[5079:5072] ,data[5087:5080] ,data[5095:5088] ,data[5287:5280] ,data[5295:5288] ,data[5303:5296] ,data[5311:5304] ,data[5319:5312] ,data[5511:5504] ,data[5519:5512] ,data[5527:5520] ,data[5535:5528] ,data[5543:5536] };
end
635 :begin
 dPIn = {data[4623:4616] ,data[4631:4624] ,data[4639:4632] ,data[4647:4640] ,data[4655:4648] ,data[4847:4840] ,data[4855:4848] ,data[4863:4856] ,data[4871:4864] ,data[4879:4872] ,data[5071:5064] ,data[5079:5072] ,data[5087:5080] ,data[5095:5088] ,data[5103:5096] ,data[5295:5288] ,data[5303:5296] ,data[5311:5304] ,data[5319:5312] ,data[5327:5320] ,data[5519:5512] ,data[5527:5520] ,data[5535:5528] ,data[5543:5536] ,data[5551:5544] };
end
636 :begin
 dPIn = {data[4631:4624] ,data[4639:4632] ,data[4647:4640] ,data[4655:4648] ,data[4663:4656] ,data[4855:4848] ,data[4863:4856] ,data[4871:4864] ,data[4879:4872] ,data[4887:4880] ,data[5079:5072] ,data[5087:5080] ,data[5095:5088] ,data[5103:5096] ,data[5111:5104] ,data[5303:5296] ,data[5311:5304] ,data[5319:5312] ,data[5327:5320] ,data[5335:5328] ,data[5527:5520] ,data[5535:5528] ,data[5543:5536] ,data[5551:5544] ,data[5559:5552] };
end
637 :begin
 dPIn = {data[4639:4632] ,data[4647:4640] ,data[4655:4648] ,data[4663:4656] ,data[4671:4664] ,data[4863:4856] ,data[4871:4864] ,data[4879:4872] ,data[4887:4880] ,data[4895:4888] ,data[5087:5080] ,data[5095:5088] ,data[5103:5096] ,data[5111:5104] ,data[5119:5112] ,data[5311:5304] ,data[5319:5312] ,data[5327:5320] ,data[5335:5328] ,data[5343:5336] ,data[5535:5528] ,data[5543:5536] ,data[5551:5544] ,data[5559:5552] ,data[5567:5560] };
end
638 :begin
 dPIn = {data[4647:4640] ,data[4655:4648] ,data[4663:4656] ,data[4671:4664] ,data[4679:4672] ,data[4871:4864] ,data[4879:4872] ,data[4887:4880] ,data[4895:4888] ,data[4903:4896] ,data[5095:5088] ,data[5103:5096] ,data[5111:5104] ,data[5119:5112] ,data[5127:5120] ,data[5319:5312] ,data[5327:5320] ,data[5335:5328] ,data[5343:5336] ,data[5351:5344] ,data[5543:5536] ,data[5551:5544] ,data[5559:5552] ,data[5567:5560] ,data[5575:5568] };
end
639 :begin
 dPIn = {data[4655:4648] ,data[4663:4656] ,data[4671:4664] ,data[4679:4672] ,data[4687:4680] ,data[4879:4872] ,data[4887:4880] ,data[4895:4888] ,data[4903:4896] ,data[4911:4904] ,data[5103:5096] ,data[5111:5104] ,data[5119:5112] ,data[5127:5120] ,data[5135:5128] ,data[5327:5320] ,data[5335:5328] ,data[5343:5336] ,data[5351:5344] ,data[5359:5352] ,data[5551:5544] ,data[5559:5552] ,data[5567:5560] ,data[5575:5568] ,data[5583:5576] };
end
640 :begin
 dPIn = {data[4663:4656] ,data[4671:4664] ,data[4679:4672] ,data[4687:4680] ,data[4695:4688] ,data[4887:4880] ,data[4895:4888] ,data[4903:4896] ,data[4911:4904] ,data[4919:4912] ,data[5111:5104] ,data[5119:5112] ,data[5127:5120] ,data[5135:5128] ,data[5143:5136] ,data[5335:5328] ,data[5343:5336] ,data[5351:5344] ,data[5359:5352] ,data[5367:5360] ,data[5559:5552] ,data[5567:5560] ,data[5575:5568] ,data[5583:5576] ,data[5591:5584] };
end
641 :begin
 dPIn = {data[4671:4664] ,data[4679:4672] ,data[4687:4680] ,data[4695:4688] ,data[4703:4696] ,data[4895:4888] ,data[4903:4896] ,data[4911:4904] ,data[4919:4912] ,data[4927:4920] ,data[5119:5112] ,data[5127:5120] ,data[5135:5128] ,data[5143:5136] ,data[5151:5144] ,data[5343:5336] ,data[5351:5344] ,data[5359:5352] ,data[5367:5360] ,data[5375:5368] ,data[5567:5560] ,data[5575:5568] ,data[5583:5576] ,data[5591:5584] ,data[5599:5592] };
end
642 :begin
 dPIn = {data[4679:4672] ,data[4687:4680] ,data[4695:4688] ,data[4703:4696] ,0 ,data[4903:4896] ,data[4911:4904] ,data[4919:4912] ,data[4927:4920] ,0 ,data[5127:5120] ,data[5135:5128] ,data[5143:5136] ,data[5151:5144] ,0 ,data[5351:5344] ,data[5359:5352] ,data[5367:5360] ,data[5375:5368] ,0 ,data[5575:5568] ,data[5583:5576] ,data[5591:5584] ,data[5599:5592] ,0 };
end
643 :begin
 dPIn = {data[4687:4680] ,data[4695:4688] ,data[4703:4696] ,0 ,0 ,data[4911:4904] ,data[4919:4912] ,data[4927:4920] ,0 ,0 ,data[5135:5128] ,data[5143:5136] ,data[5151:5144] ,0 ,0 ,data[5359:5352] ,data[5367:5360] ,data[5375:5368] ,0 ,0 ,data[5583:5576] ,data[5591:5584] ,data[5599:5592] ,0 ,0 };
end
644 :begin
 dPIn = {0 ,0 ,data[4711:4704] ,data[4719:4712] ,data[4727:4720] ,0 ,0 ,data[4935:4928] ,data[4943:4936] ,data[4951:4944] ,0 ,0 ,data[5159:5152] ,data[5167:5160] ,data[5175:5168] ,0 ,0 ,data[5383:5376] ,data[5391:5384] ,data[5399:5392] ,0 ,0 ,data[5607:5600] ,data[5615:5608] ,data[5623:5616] };
end
645 :begin
 dPIn = {0 ,data[4711:4704] ,data[4719:4712] ,data[4727:4720] ,data[4735:4728] ,0 ,data[4935:4928] ,data[4943:4936] ,data[4951:4944] ,data[4959:4952] ,0 ,data[5159:5152] ,data[5167:5160] ,data[5175:5168] ,data[5183:5176] ,0 ,data[5383:5376] ,data[5391:5384] ,data[5399:5392] ,data[5407:5400] ,0 ,data[5607:5600] ,data[5615:5608] ,data[5623:5616] ,data[5631:5624] };
end
646 :begin
 dPIn = {data[4711:4704] ,data[4719:4712] ,data[4727:4720] ,data[4735:4728] ,data[4743:4736] ,data[4935:4928] ,data[4943:4936] ,data[4951:4944] ,data[4959:4952] ,data[4967:4960] ,data[5159:5152] ,data[5167:5160] ,data[5175:5168] ,data[5183:5176] ,data[5191:5184] ,data[5383:5376] ,data[5391:5384] ,data[5399:5392] ,data[5407:5400] ,data[5415:5408] ,data[5607:5600] ,data[5615:5608] ,data[5623:5616] ,data[5631:5624] ,data[5639:5632] };
end
647 :begin
 dPIn = {data[4719:4712] ,data[4727:4720] ,data[4735:4728] ,data[4743:4736] ,data[4751:4744] ,data[4943:4936] ,data[4951:4944] ,data[4959:4952] ,data[4967:4960] ,data[4975:4968] ,data[5167:5160] ,data[5175:5168] ,data[5183:5176] ,data[5191:5184] ,data[5199:5192] ,data[5391:5384] ,data[5399:5392] ,data[5407:5400] ,data[5415:5408] ,data[5423:5416] ,data[5615:5608] ,data[5623:5616] ,data[5631:5624] ,data[5639:5632] ,data[5647:5640] };
end
648 :begin
 dPIn = {data[4727:4720] ,data[4735:4728] ,data[4743:4736] ,data[4751:4744] ,data[4759:4752] ,data[4951:4944] ,data[4959:4952] ,data[4967:4960] ,data[4975:4968] ,data[4983:4976] ,data[5175:5168] ,data[5183:5176] ,data[5191:5184] ,data[5199:5192] ,data[5207:5200] ,data[5399:5392] ,data[5407:5400] ,data[5415:5408] ,data[5423:5416] ,data[5431:5424] ,data[5623:5616] ,data[5631:5624] ,data[5639:5632] ,data[5647:5640] ,data[5655:5648] };
end
649 :begin
 dPIn = {data[4735:4728] ,data[4743:4736] ,data[4751:4744] ,data[4759:4752] ,data[4767:4760] ,data[4959:4952] ,data[4967:4960] ,data[4975:4968] ,data[4983:4976] ,data[4991:4984] ,data[5183:5176] ,data[5191:5184] ,data[5199:5192] ,data[5207:5200] ,data[5215:5208] ,data[5407:5400] ,data[5415:5408] ,data[5423:5416] ,data[5431:5424] ,data[5439:5432] ,data[5631:5624] ,data[5639:5632] ,data[5647:5640] ,data[5655:5648] ,data[5663:5656] };
end
650 :begin
 dPIn = {data[4743:4736] ,data[4751:4744] ,data[4759:4752] ,data[4767:4760] ,data[4775:4768] ,data[4967:4960] ,data[4975:4968] ,data[4983:4976] ,data[4991:4984] ,data[4999:4992] ,data[5191:5184] ,data[5199:5192] ,data[5207:5200] ,data[5215:5208] ,data[5223:5216] ,data[5415:5408] ,data[5423:5416] ,data[5431:5424] ,data[5439:5432] ,data[5447:5440] ,data[5639:5632] ,data[5647:5640] ,data[5655:5648] ,data[5663:5656] ,data[5671:5664] };
end
651 :begin
 dPIn = {data[4751:4744] ,data[4759:4752] ,data[4767:4760] ,data[4775:4768] ,data[4783:4776] ,data[4975:4968] ,data[4983:4976] ,data[4991:4984] ,data[4999:4992] ,data[5007:5000] ,data[5199:5192] ,data[5207:5200] ,data[5215:5208] ,data[5223:5216] ,data[5231:5224] ,data[5423:5416] ,data[5431:5424] ,data[5439:5432] ,data[5447:5440] ,data[5455:5448] ,data[5647:5640] ,data[5655:5648] ,data[5663:5656] ,data[5671:5664] ,data[5679:5672] };
end
652 :begin
 dPIn = {data[4759:4752] ,data[4767:4760] ,data[4775:4768] ,data[4783:4776] ,data[4791:4784] ,data[4983:4976] ,data[4991:4984] ,data[4999:4992] ,data[5007:5000] ,data[5015:5008] ,data[5207:5200] ,data[5215:5208] ,data[5223:5216] ,data[5231:5224] ,data[5239:5232] ,data[5431:5424] ,data[5439:5432] ,data[5447:5440] ,data[5455:5448] ,data[5463:5456] ,data[5655:5648] ,data[5663:5656] ,data[5671:5664] ,data[5679:5672] ,data[5687:5680] };
end
653 :begin
 dPIn = {data[4767:4760] ,data[4775:4768] ,data[4783:4776] ,data[4791:4784] ,data[4799:4792] ,data[4991:4984] ,data[4999:4992] ,data[5007:5000] ,data[5015:5008] ,data[5023:5016] ,data[5215:5208] ,data[5223:5216] ,data[5231:5224] ,data[5239:5232] ,data[5247:5240] ,data[5439:5432] ,data[5447:5440] ,data[5455:5448] ,data[5463:5456] ,data[5471:5464] ,data[5663:5656] ,data[5671:5664] ,data[5679:5672] ,data[5687:5680] ,data[5695:5688] };
end
654 :begin
 dPIn = {data[4775:4768] ,data[4783:4776] ,data[4791:4784] ,data[4799:4792] ,data[4807:4800] ,data[4999:4992] ,data[5007:5000] ,data[5015:5008] ,data[5023:5016] ,data[5031:5024] ,data[5223:5216] ,data[5231:5224] ,data[5239:5232] ,data[5247:5240] ,data[5255:5248] ,data[5447:5440] ,data[5455:5448] ,data[5463:5456] ,data[5471:5464] ,data[5479:5472] ,data[5671:5664] ,data[5679:5672] ,data[5687:5680] ,data[5695:5688] ,data[5703:5696] };
end
655 :begin
 dPIn = {data[4783:4776] ,data[4791:4784] ,data[4799:4792] ,data[4807:4800] ,data[4815:4808] ,data[5007:5000] ,data[5015:5008] ,data[5023:5016] ,data[5031:5024] ,data[5039:5032] ,data[5231:5224] ,data[5239:5232] ,data[5247:5240] ,data[5255:5248] ,data[5263:5256] ,data[5455:5448] ,data[5463:5456] ,data[5471:5464] ,data[5479:5472] ,data[5487:5480] ,data[5679:5672] ,data[5687:5680] ,data[5695:5688] ,data[5703:5696] ,data[5711:5704] };
end
656 :begin
 dPIn = {data[4791:4784] ,data[4799:4792] ,data[4807:4800] ,data[4815:4808] ,data[4823:4816] ,data[5015:5008] ,data[5023:5016] ,data[5031:5024] ,data[5039:5032] ,data[5047:5040] ,data[5239:5232] ,data[5247:5240] ,data[5255:5248] ,data[5263:5256] ,data[5271:5264] ,data[5463:5456] ,data[5471:5464] ,data[5479:5472] ,data[5487:5480] ,data[5495:5488] ,data[5687:5680] ,data[5695:5688] ,data[5703:5696] ,data[5711:5704] ,data[5719:5712] };
end
657 :begin
 dPIn = {data[4799:4792] ,data[4807:4800] ,data[4815:4808] ,data[4823:4816] ,data[4831:4824] ,data[5023:5016] ,data[5031:5024] ,data[5039:5032] ,data[5047:5040] ,data[5055:5048] ,data[5247:5240] ,data[5255:5248] ,data[5263:5256] ,data[5271:5264] ,data[5279:5272] ,data[5471:5464] ,data[5479:5472] ,data[5487:5480] ,data[5495:5488] ,data[5503:5496] ,data[5695:5688] ,data[5703:5696] ,data[5711:5704] ,data[5719:5712] ,data[5727:5720] };
end
658 :begin
 dPIn = {data[4807:4800] ,data[4815:4808] ,data[4823:4816] ,data[4831:4824] ,data[4839:4832] ,data[5031:5024] ,data[5039:5032] ,data[5047:5040] ,data[5055:5048] ,data[5063:5056] ,data[5255:5248] ,data[5263:5256] ,data[5271:5264] ,data[5279:5272] ,data[5287:5280] ,data[5479:5472] ,data[5487:5480] ,data[5495:5488] ,data[5503:5496] ,data[5511:5504] ,data[5703:5696] ,data[5711:5704] ,data[5719:5712] ,data[5727:5720] ,data[5735:5728] };
end
659 :begin
 dPIn = {data[4815:4808] ,data[4823:4816] ,data[4831:4824] ,data[4839:4832] ,data[4847:4840] ,data[5039:5032] ,data[5047:5040] ,data[5055:5048] ,data[5063:5056] ,data[5071:5064] ,data[5263:5256] ,data[5271:5264] ,data[5279:5272] ,data[5287:5280] ,data[5295:5288] ,data[5487:5480] ,data[5495:5488] ,data[5503:5496] ,data[5511:5504] ,data[5519:5512] ,data[5711:5704] ,data[5719:5712] ,data[5727:5720] ,data[5735:5728] ,data[5743:5736] };
end
660 :begin
 dPIn = {data[4823:4816] ,data[4831:4824] ,data[4839:4832] ,data[4847:4840] ,data[4855:4848] ,data[5047:5040] ,data[5055:5048] ,data[5063:5056] ,data[5071:5064] ,data[5079:5072] ,data[5271:5264] ,data[5279:5272] ,data[5287:5280] ,data[5295:5288] ,data[5303:5296] ,data[5495:5488] ,data[5503:5496] ,data[5511:5504] ,data[5519:5512] ,data[5527:5520] ,data[5719:5712] ,data[5727:5720] ,data[5735:5728] ,data[5743:5736] ,data[5751:5744] };
end
661 :begin
 dPIn = {data[4831:4824] ,data[4839:4832] ,data[4847:4840] ,data[4855:4848] ,data[4863:4856] ,data[5055:5048] ,data[5063:5056] ,data[5071:5064] ,data[5079:5072] ,data[5087:5080] ,data[5279:5272] ,data[5287:5280] ,data[5295:5288] ,data[5303:5296] ,data[5311:5304] ,data[5503:5496] ,data[5511:5504] ,data[5519:5512] ,data[5527:5520] ,data[5535:5528] ,data[5727:5720] ,data[5735:5728] ,data[5743:5736] ,data[5751:5744] ,data[5759:5752] };
end
662 :begin
 dPIn = {data[4839:4832] ,data[4847:4840] ,data[4855:4848] ,data[4863:4856] ,data[4871:4864] ,data[5063:5056] ,data[5071:5064] ,data[5079:5072] ,data[5087:5080] ,data[5095:5088] ,data[5287:5280] ,data[5295:5288] ,data[5303:5296] ,data[5311:5304] ,data[5319:5312] ,data[5511:5504] ,data[5519:5512] ,data[5527:5520] ,data[5535:5528] ,data[5543:5536] ,data[5735:5728] ,data[5743:5736] ,data[5751:5744] ,data[5759:5752] ,data[5767:5760] };
end
663 :begin
 dPIn = {data[4847:4840] ,data[4855:4848] ,data[4863:4856] ,data[4871:4864] ,data[4879:4872] ,data[5071:5064] ,data[5079:5072] ,data[5087:5080] ,data[5095:5088] ,data[5103:5096] ,data[5295:5288] ,data[5303:5296] ,data[5311:5304] ,data[5319:5312] ,data[5327:5320] ,data[5519:5512] ,data[5527:5520] ,data[5535:5528] ,data[5543:5536] ,data[5551:5544] ,data[5743:5736] ,data[5751:5744] ,data[5759:5752] ,data[5767:5760] ,data[5775:5768] };
end
664 :begin
 dPIn = {data[4855:4848] ,data[4863:4856] ,data[4871:4864] ,data[4879:4872] ,data[4887:4880] ,data[5079:5072] ,data[5087:5080] ,data[5095:5088] ,data[5103:5096] ,data[5111:5104] ,data[5303:5296] ,data[5311:5304] ,data[5319:5312] ,data[5327:5320] ,data[5335:5328] ,data[5527:5520] ,data[5535:5528] ,data[5543:5536] ,data[5551:5544] ,data[5559:5552] ,data[5751:5744] ,data[5759:5752] ,data[5767:5760] ,data[5775:5768] ,data[5783:5776] };
end
665 :begin
 dPIn = {data[4863:4856] ,data[4871:4864] ,data[4879:4872] ,data[4887:4880] ,data[4895:4888] ,data[5087:5080] ,data[5095:5088] ,data[5103:5096] ,data[5111:5104] ,data[5119:5112] ,data[5311:5304] ,data[5319:5312] ,data[5327:5320] ,data[5335:5328] ,data[5343:5336] ,data[5535:5528] ,data[5543:5536] ,data[5551:5544] ,data[5559:5552] ,data[5567:5560] ,data[5759:5752] ,data[5767:5760] ,data[5775:5768] ,data[5783:5776] ,data[5791:5784] };
end
666 :begin
 dPIn = {data[4871:4864] ,data[4879:4872] ,data[4887:4880] ,data[4895:4888] ,data[4903:4896] ,data[5095:5088] ,data[5103:5096] ,data[5111:5104] ,data[5119:5112] ,data[5127:5120] ,data[5319:5312] ,data[5327:5320] ,data[5335:5328] ,data[5343:5336] ,data[5351:5344] ,data[5543:5536] ,data[5551:5544] ,data[5559:5552] ,data[5567:5560] ,data[5575:5568] ,data[5767:5760] ,data[5775:5768] ,data[5783:5776] ,data[5791:5784] ,data[5799:5792] };
end
667 :begin
 dPIn = {data[4879:4872] ,data[4887:4880] ,data[4895:4888] ,data[4903:4896] ,data[4911:4904] ,data[5103:5096] ,data[5111:5104] ,data[5119:5112] ,data[5127:5120] ,data[5135:5128] ,data[5327:5320] ,data[5335:5328] ,data[5343:5336] ,data[5351:5344] ,data[5359:5352] ,data[5551:5544] ,data[5559:5552] ,data[5567:5560] ,data[5575:5568] ,data[5583:5576] ,data[5775:5768] ,data[5783:5776] ,data[5791:5784] ,data[5799:5792] ,data[5807:5800] };
end
668 :begin
 dPIn = {data[4887:4880] ,data[4895:4888] ,data[4903:4896] ,data[4911:4904] ,data[4919:4912] ,data[5111:5104] ,data[5119:5112] ,data[5127:5120] ,data[5135:5128] ,data[5143:5136] ,data[5335:5328] ,data[5343:5336] ,data[5351:5344] ,data[5359:5352] ,data[5367:5360] ,data[5559:5552] ,data[5567:5560] ,data[5575:5568] ,data[5583:5576] ,data[5591:5584] ,data[5783:5776] ,data[5791:5784] ,data[5799:5792] ,data[5807:5800] ,data[5815:5808] };
end
669 :begin
 dPIn = {data[4895:4888] ,data[4903:4896] ,data[4911:4904] ,data[4919:4912] ,data[4927:4920] ,data[5119:5112] ,data[5127:5120] ,data[5135:5128] ,data[5143:5136] ,data[5151:5144] ,data[5343:5336] ,data[5351:5344] ,data[5359:5352] ,data[5367:5360] ,data[5375:5368] ,data[5567:5560] ,data[5575:5568] ,data[5583:5576] ,data[5591:5584] ,data[5599:5592] ,data[5791:5784] ,data[5799:5792] ,data[5807:5800] ,data[5815:5808] ,data[5823:5816] };
end
670 :begin
 dPIn = {data[4903:4896] ,data[4911:4904] ,data[4919:4912] ,data[4927:4920] ,0 ,data[5127:5120] ,data[5135:5128] ,data[5143:5136] ,data[5151:5144] ,0 ,data[5351:5344] ,data[5359:5352] ,data[5367:5360] ,data[5375:5368] ,0 ,data[5575:5568] ,data[5583:5576] ,data[5591:5584] ,data[5599:5592] ,0 ,data[5799:5792] ,data[5807:5800] ,data[5815:5808] ,data[5823:5816] ,0 };
end
671 :begin
 dPIn = {data[4911:4904] ,data[4919:4912] ,data[4927:4920] ,0 ,0 ,data[5135:5128] ,data[5143:5136] ,data[5151:5144] ,0 ,0 ,data[5359:5352] ,data[5367:5360] ,data[5375:5368] ,0 ,0 ,data[5583:5576] ,data[5591:5584] ,data[5599:5592] ,0 ,0 ,data[5807:5800] ,data[5815:5808] ,data[5823:5816] ,0 ,0 };
end
672 :begin
 dPIn = {0 ,0 ,data[4935:4928] ,data[4943:4936] ,data[4951:4944] ,0 ,0 ,data[5159:5152] ,data[5167:5160] ,data[5175:5168] ,0 ,0 ,data[5383:5376] ,data[5391:5384] ,data[5399:5392] ,0 ,0 ,data[5607:5600] ,data[5615:5608] ,data[5623:5616] ,0 ,0 ,data[5831:5824] ,data[5839:5832] ,data[5847:5840] };
end
673 :begin
 dPIn = {0 ,data[4935:4928] ,data[4943:4936] ,data[4951:4944] ,data[4959:4952] ,0 ,data[5159:5152] ,data[5167:5160] ,data[5175:5168] ,data[5183:5176] ,0 ,data[5383:5376] ,data[5391:5384] ,data[5399:5392] ,data[5407:5400] ,0 ,data[5607:5600] ,data[5615:5608] ,data[5623:5616] ,data[5631:5624] ,0 ,data[5831:5824] ,data[5839:5832] ,data[5847:5840] ,data[5855:5848] };
end
674 :begin
 dPIn = {data[4935:4928] ,data[4943:4936] ,data[4951:4944] ,data[4959:4952] ,data[4967:4960] ,data[5159:5152] ,data[5167:5160] ,data[5175:5168] ,data[5183:5176] ,data[5191:5184] ,data[5383:5376] ,data[5391:5384] ,data[5399:5392] ,data[5407:5400] ,data[5415:5408] ,data[5607:5600] ,data[5615:5608] ,data[5623:5616] ,data[5631:5624] ,data[5639:5632] ,data[5831:5824] ,data[5839:5832] ,data[5847:5840] ,data[5855:5848] ,data[5863:5856] };
end
675 :begin
 dPIn = {data[4943:4936] ,data[4951:4944] ,data[4959:4952] ,data[4967:4960] ,data[4975:4968] ,data[5167:5160] ,data[5175:5168] ,data[5183:5176] ,data[5191:5184] ,data[5199:5192] ,data[5391:5384] ,data[5399:5392] ,data[5407:5400] ,data[5415:5408] ,data[5423:5416] ,data[5615:5608] ,data[5623:5616] ,data[5631:5624] ,data[5639:5632] ,data[5647:5640] ,data[5839:5832] ,data[5847:5840] ,data[5855:5848] ,data[5863:5856] ,data[5871:5864] };
end
676 :begin
 dPIn = {data[4951:4944] ,data[4959:4952] ,data[4967:4960] ,data[4975:4968] ,data[4983:4976] ,data[5175:5168] ,data[5183:5176] ,data[5191:5184] ,data[5199:5192] ,data[5207:5200] ,data[5399:5392] ,data[5407:5400] ,data[5415:5408] ,data[5423:5416] ,data[5431:5424] ,data[5623:5616] ,data[5631:5624] ,data[5639:5632] ,data[5647:5640] ,data[5655:5648] ,data[5847:5840] ,data[5855:5848] ,data[5863:5856] ,data[5871:5864] ,data[5879:5872] };
end
677 :begin
 dPIn = {data[4959:4952] ,data[4967:4960] ,data[4975:4968] ,data[4983:4976] ,data[4991:4984] ,data[5183:5176] ,data[5191:5184] ,data[5199:5192] ,data[5207:5200] ,data[5215:5208] ,data[5407:5400] ,data[5415:5408] ,data[5423:5416] ,data[5431:5424] ,data[5439:5432] ,data[5631:5624] ,data[5639:5632] ,data[5647:5640] ,data[5655:5648] ,data[5663:5656] ,data[5855:5848] ,data[5863:5856] ,data[5871:5864] ,data[5879:5872] ,data[5887:5880] };
end
678 :begin
 dPIn = {data[4967:4960] ,data[4975:4968] ,data[4983:4976] ,data[4991:4984] ,data[4999:4992] ,data[5191:5184] ,data[5199:5192] ,data[5207:5200] ,data[5215:5208] ,data[5223:5216] ,data[5415:5408] ,data[5423:5416] ,data[5431:5424] ,data[5439:5432] ,data[5447:5440] ,data[5639:5632] ,data[5647:5640] ,data[5655:5648] ,data[5663:5656] ,data[5671:5664] ,data[5863:5856] ,data[5871:5864] ,data[5879:5872] ,data[5887:5880] ,data[5895:5888] };
end
679 :begin
 dPIn = {data[4975:4968] ,data[4983:4976] ,data[4991:4984] ,data[4999:4992] ,data[5007:5000] ,data[5199:5192] ,data[5207:5200] ,data[5215:5208] ,data[5223:5216] ,data[5231:5224] ,data[5423:5416] ,data[5431:5424] ,data[5439:5432] ,data[5447:5440] ,data[5455:5448] ,data[5647:5640] ,data[5655:5648] ,data[5663:5656] ,data[5671:5664] ,data[5679:5672] ,data[5871:5864] ,data[5879:5872] ,data[5887:5880] ,data[5895:5888] ,data[5903:5896] };
end
680 :begin
 dPIn = {data[4983:4976] ,data[4991:4984] ,data[4999:4992] ,data[5007:5000] ,data[5015:5008] ,data[5207:5200] ,data[5215:5208] ,data[5223:5216] ,data[5231:5224] ,data[5239:5232] ,data[5431:5424] ,data[5439:5432] ,data[5447:5440] ,data[5455:5448] ,data[5463:5456] ,data[5655:5648] ,data[5663:5656] ,data[5671:5664] ,data[5679:5672] ,data[5687:5680] ,data[5879:5872] ,data[5887:5880] ,data[5895:5888] ,data[5903:5896] ,data[5911:5904] };
end
681 :begin
 dPIn = {data[4991:4984] ,data[4999:4992] ,data[5007:5000] ,data[5015:5008] ,data[5023:5016] ,data[5215:5208] ,data[5223:5216] ,data[5231:5224] ,data[5239:5232] ,data[5247:5240] ,data[5439:5432] ,data[5447:5440] ,data[5455:5448] ,data[5463:5456] ,data[5471:5464] ,data[5663:5656] ,data[5671:5664] ,data[5679:5672] ,data[5687:5680] ,data[5695:5688] ,data[5887:5880] ,data[5895:5888] ,data[5903:5896] ,data[5911:5904] ,data[5919:5912] };
end
682 :begin
 dPIn = {data[4999:4992] ,data[5007:5000] ,data[5015:5008] ,data[5023:5016] ,data[5031:5024] ,data[5223:5216] ,data[5231:5224] ,data[5239:5232] ,data[5247:5240] ,data[5255:5248] ,data[5447:5440] ,data[5455:5448] ,data[5463:5456] ,data[5471:5464] ,data[5479:5472] ,data[5671:5664] ,data[5679:5672] ,data[5687:5680] ,data[5695:5688] ,data[5703:5696] ,data[5895:5888] ,data[5903:5896] ,data[5911:5904] ,data[5919:5912] ,data[5927:5920] };
end
683 :begin
 dPIn = {data[5007:5000] ,data[5015:5008] ,data[5023:5016] ,data[5031:5024] ,data[5039:5032] ,data[5231:5224] ,data[5239:5232] ,data[5247:5240] ,data[5255:5248] ,data[5263:5256] ,data[5455:5448] ,data[5463:5456] ,data[5471:5464] ,data[5479:5472] ,data[5487:5480] ,data[5679:5672] ,data[5687:5680] ,data[5695:5688] ,data[5703:5696] ,data[5711:5704] ,data[5903:5896] ,data[5911:5904] ,data[5919:5912] ,data[5927:5920] ,data[5935:5928] };
end
684 :begin
 dPIn = {data[5015:5008] ,data[5023:5016] ,data[5031:5024] ,data[5039:5032] ,data[5047:5040] ,data[5239:5232] ,data[5247:5240] ,data[5255:5248] ,data[5263:5256] ,data[5271:5264] ,data[5463:5456] ,data[5471:5464] ,data[5479:5472] ,data[5487:5480] ,data[5495:5488] ,data[5687:5680] ,data[5695:5688] ,data[5703:5696] ,data[5711:5704] ,data[5719:5712] ,data[5911:5904] ,data[5919:5912] ,data[5927:5920] ,data[5935:5928] ,data[5943:5936] };
end
685 :begin
 dPIn = {data[5023:5016] ,data[5031:5024] ,data[5039:5032] ,data[5047:5040] ,data[5055:5048] ,data[5247:5240] ,data[5255:5248] ,data[5263:5256] ,data[5271:5264] ,data[5279:5272] ,data[5471:5464] ,data[5479:5472] ,data[5487:5480] ,data[5495:5488] ,data[5503:5496] ,data[5695:5688] ,data[5703:5696] ,data[5711:5704] ,data[5719:5712] ,data[5727:5720] ,data[5919:5912] ,data[5927:5920] ,data[5935:5928] ,data[5943:5936] ,data[5951:5944] };
end
686 :begin
 dPIn = {data[5031:5024] ,data[5039:5032] ,data[5047:5040] ,data[5055:5048] ,data[5063:5056] ,data[5255:5248] ,data[5263:5256] ,data[5271:5264] ,data[5279:5272] ,data[5287:5280] ,data[5479:5472] ,data[5487:5480] ,data[5495:5488] ,data[5503:5496] ,data[5511:5504] ,data[5703:5696] ,data[5711:5704] ,data[5719:5712] ,data[5727:5720] ,data[5735:5728] ,data[5927:5920] ,data[5935:5928] ,data[5943:5936] ,data[5951:5944] ,data[5959:5952] };
end
687 :begin
 dPIn = {data[5039:5032] ,data[5047:5040] ,data[5055:5048] ,data[5063:5056] ,data[5071:5064] ,data[5263:5256] ,data[5271:5264] ,data[5279:5272] ,data[5287:5280] ,data[5295:5288] ,data[5487:5480] ,data[5495:5488] ,data[5503:5496] ,data[5511:5504] ,data[5519:5512] ,data[5711:5704] ,data[5719:5712] ,data[5727:5720] ,data[5735:5728] ,data[5743:5736] ,data[5935:5928] ,data[5943:5936] ,data[5951:5944] ,data[5959:5952] ,data[5967:5960] };
end
688 :begin
 dPIn = {data[5047:5040] ,data[5055:5048] ,data[5063:5056] ,data[5071:5064] ,data[5079:5072] ,data[5271:5264] ,data[5279:5272] ,data[5287:5280] ,data[5295:5288] ,data[5303:5296] ,data[5495:5488] ,data[5503:5496] ,data[5511:5504] ,data[5519:5512] ,data[5527:5520] ,data[5719:5712] ,data[5727:5720] ,data[5735:5728] ,data[5743:5736] ,data[5751:5744] ,data[5943:5936] ,data[5951:5944] ,data[5959:5952] ,data[5967:5960] ,data[5975:5968] };
end
689 :begin
 dPIn = {data[5055:5048] ,data[5063:5056] ,data[5071:5064] ,data[5079:5072] ,data[5087:5080] ,data[5279:5272] ,data[5287:5280] ,data[5295:5288] ,data[5303:5296] ,data[5311:5304] ,data[5503:5496] ,data[5511:5504] ,data[5519:5512] ,data[5527:5520] ,data[5535:5528] ,data[5727:5720] ,data[5735:5728] ,data[5743:5736] ,data[5751:5744] ,data[5759:5752] ,data[5951:5944] ,data[5959:5952] ,data[5967:5960] ,data[5975:5968] ,data[5983:5976] };
end
690 :begin
 dPIn = {data[5063:5056] ,data[5071:5064] ,data[5079:5072] ,data[5087:5080] ,data[5095:5088] ,data[5287:5280] ,data[5295:5288] ,data[5303:5296] ,data[5311:5304] ,data[5319:5312] ,data[5511:5504] ,data[5519:5512] ,data[5527:5520] ,data[5535:5528] ,data[5543:5536] ,data[5735:5728] ,data[5743:5736] ,data[5751:5744] ,data[5759:5752] ,data[5767:5760] ,data[5959:5952] ,data[5967:5960] ,data[5975:5968] ,data[5983:5976] ,data[5991:5984] };
end
691 :begin
 dPIn = {data[5071:5064] ,data[5079:5072] ,data[5087:5080] ,data[5095:5088] ,data[5103:5096] ,data[5295:5288] ,data[5303:5296] ,data[5311:5304] ,data[5319:5312] ,data[5327:5320] ,data[5519:5512] ,data[5527:5520] ,data[5535:5528] ,data[5543:5536] ,data[5551:5544] ,data[5743:5736] ,data[5751:5744] ,data[5759:5752] ,data[5767:5760] ,data[5775:5768] ,data[5967:5960] ,data[5975:5968] ,data[5983:5976] ,data[5991:5984] ,data[5999:5992] };
end
692 :begin
 dPIn = {data[5079:5072] ,data[5087:5080] ,data[5095:5088] ,data[5103:5096] ,data[5111:5104] ,data[5303:5296] ,data[5311:5304] ,data[5319:5312] ,data[5327:5320] ,data[5335:5328] ,data[5527:5520] ,data[5535:5528] ,data[5543:5536] ,data[5551:5544] ,data[5559:5552] ,data[5751:5744] ,data[5759:5752] ,data[5767:5760] ,data[5775:5768] ,data[5783:5776] ,data[5975:5968] ,data[5983:5976] ,data[5991:5984] ,data[5999:5992] ,data[6007:6000] };
end
693 :begin
 dPIn = {data[5087:5080] ,data[5095:5088] ,data[5103:5096] ,data[5111:5104] ,data[5119:5112] ,data[5311:5304] ,data[5319:5312] ,data[5327:5320] ,data[5335:5328] ,data[5343:5336] ,data[5535:5528] ,data[5543:5536] ,data[5551:5544] ,data[5559:5552] ,data[5567:5560] ,data[5759:5752] ,data[5767:5760] ,data[5775:5768] ,data[5783:5776] ,data[5791:5784] ,data[5983:5976] ,data[5991:5984] ,data[5999:5992] ,data[6007:6000] ,data[6015:6008] };
end
694 :begin
 dPIn = {data[5095:5088] ,data[5103:5096] ,data[5111:5104] ,data[5119:5112] ,data[5127:5120] ,data[5319:5312] ,data[5327:5320] ,data[5335:5328] ,data[5343:5336] ,data[5351:5344] ,data[5543:5536] ,data[5551:5544] ,data[5559:5552] ,data[5567:5560] ,data[5575:5568] ,data[5767:5760] ,data[5775:5768] ,data[5783:5776] ,data[5791:5784] ,data[5799:5792] ,data[5991:5984] ,data[5999:5992] ,data[6007:6000] ,data[6015:6008] ,data[6023:6016] };
end
695 :begin
 dPIn = {data[5103:5096] ,data[5111:5104] ,data[5119:5112] ,data[5127:5120] ,data[5135:5128] ,data[5327:5320] ,data[5335:5328] ,data[5343:5336] ,data[5351:5344] ,data[5359:5352] ,data[5551:5544] ,data[5559:5552] ,data[5567:5560] ,data[5575:5568] ,data[5583:5576] ,data[5775:5768] ,data[5783:5776] ,data[5791:5784] ,data[5799:5792] ,data[5807:5800] ,data[5999:5992] ,data[6007:6000] ,data[6015:6008] ,data[6023:6016] ,data[6031:6024] };
end
696 :begin
 dPIn = {data[5111:5104] ,data[5119:5112] ,data[5127:5120] ,data[5135:5128] ,data[5143:5136] ,data[5335:5328] ,data[5343:5336] ,data[5351:5344] ,data[5359:5352] ,data[5367:5360] ,data[5559:5552] ,data[5567:5560] ,data[5575:5568] ,data[5583:5576] ,data[5591:5584] ,data[5783:5776] ,data[5791:5784] ,data[5799:5792] ,data[5807:5800] ,data[5815:5808] ,data[6007:6000] ,data[6015:6008] ,data[6023:6016] ,data[6031:6024] ,data[6039:6032] };
end
697 :begin
 dPIn = {data[5119:5112] ,data[5127:5120] ,data[5135:5128] ,data[5143:5136] ,data[5151:5144] ,data[5343:5336] ,data[5351:5344] ,data[5359:5352] ,data[5367:5360] ,data[5375:5368] ,data[5567:5560] ,data[5575:5568] ,data[5583:5576] ,data[5591:5584] ,data[5599:5592] ,data[5791:5784] ,data[5799:5792] ,data[5807:5800] ,data[5815:5808] ,data[5823:5816] ,data[6015:6008] ,data[6023:6016] ,data[6031:6024] ,data[6039:6032] ,data[6047:6040] };
end
698 :begin
 dPIn = {data[5127:5120] ,data[5135:5128] ,data[5143:5136] ,data[5151:5144] ,0 ,data[5351:5344] ,data[5359:5352] ,data[5367:5360] ,data[5375:5368] ,0 ,data[5575:5568] ,data[5583:5576] ,data[5591:5584] ,data[5599:5592] ,0 ,data[5799:5792] ,data[5807:5800] ,data[5815:5808] ,data[5823:5816] ,0 ,data[6023:6016] ,data[6031:6024] ,data[6039:6032] ,data[6047:6040] ,0 };
end
699 :begin
 dPIn = {data[5135:5128] ,data[5143:5136] ,data[5151:5144] ,0 ,0 ,data[5359:5352] ,data[5367:5360] ,data[5375:5368] ,0 ,0 ,data[5583:5576] ,data[5591:5584] ,data[5599:5592] ,0 ,0 ,data[5807:5800] ,data[5815:5808] ,data[5823:5816] ,0 ,0 ,data[6031:6024] ,data[6039:6032] ,data[6047:6040] ,0 ,0 };
end
700 :begin
 dPIn = {0 ,0 ,data[5159:5152] ,data[5167:5160] ,data[5175:5168] ,0 ,0 ,data[5383:5376] ,data[5391:5384] ,data[5399:5392] ,0 ,0 ,data[5607:5600] ,data[5615:5608] ,data[5623:5616] ,0 ,0 ,data[5831:5824] ,data[5839:5832] ,data[5847:5840] ,0 ,0 ,data[6055:6048] ,data[6063:6056] ,data[6071:6064] };
end
701 :begin
 dPIn = {0 ,data[5159:5152] ,data[5167:5160] ,data[5175:5168] ,data[5183:5176] ,0 ,data[5383:5376] ,data[5391:5384] ,data[5399:5392] ,data[5407:5400] ,0 ,data[5607:5600] ,data[5615:5608] ,data[5623:5616] ,data[5631:5624] ,0 ,data[5831:5824] ,data[5839:5832] ,data[5847:5840] ,data[5855:5848] ,0 ,data[6055:6048] ,data[6063:6056] ,data[6071:6064] ,data[6079:6072] };
end
702 :begin
 dPIn = {data[5159:5152] ,data[5167:5160] ,data[5175:5168] ,data[5183:5176] ,data[5191:5184] ,data[5383:5376] ,data[5391:5384] ,data[5399:5392] ,data[5407:5400] ,data[5415:5408] ,data[5607:5600] ,data[5615:5608] ,data[5623:5616] ,data[5631:5624] ,data[5639:5632] ,data[5831:5824] ,data[5839:5832] ,data[5847:5840] ,data[5855:5848] ,data[5863:5856] ,data[6055:6048] ,data[6063:6056] ,data[6071:6064] ,data[6079:6072] ,data[6087:6080] };
end
703 :begin
 dPIn = {data[5167:5160] ,data[5175:5168] ,data[5183:5176] ,data[5191:5184] ,data[5199:5192] ,data[5391:5384] ,data[5399:5392] ,data[5407:5400] ,data[5415:5408] ,data[5423:5416] ,data[5615:5608] ,data[5623:5616] ,data[5631:5624] ,data[5639:5632] ,data[5647:5640] ,data[5839:5832] ,data[5847:5840] ,data[5855:5848] ,data[5863:5856] ,data[5871:5864] ,data[6063:6056] ,data[6071:6064] ,data[6079:6072] ,data[6087:6080] ,data[6095:6088] };
end
704 :begin
 dPIn = {data[5175:5168] ,data[5183:5176] ,data[5191:5184] ,data[5199:5192] ,data[5207:5200] ,data[5399:5392] ,data[5407:5400] ,data[5415:5408] ,data[5423:5416] ,data[5431:5424] ,data[5623:5616] ,data[5631:5624] ,data[5639:5632] ,data[5647:5640] ,data[5655:5648] ,data[5847:5840] ,data[5855:5848] ,data[5863:5856] ,data[5871:5864] ,data[5879:5872] ,data[6071:6064] ,data[6079:6072] ,data[6087:6080] ,data[6095:6088] ,data[6103:6096] };
end
705 :begin
 dPIn = {data[5183:5176] ,data[5191:5184] ,data[5199:5192] ,data[5207:5200] ,data[5215:5208] ,data[5407:5400] ,data[5415:5408] ,data[5423:5416] ,data[5431:5424] ,data[5439:5432] ,data[5631:5624] ,data[5639:5632] ,data[5647:5640] ,data[5655:5648] ,data[5663:5656] ,data[5855:5848] ,data[5863:5856] ,data[5871:5864] ,data[5879:5872] ,data[5887:5880] ,data[6079:6072] ,data[6087:6080] ,data[6095:6088] ,data[6103:6096] ,data[6111:6104] };
end
706 :begin
 dPIn = {data[5191:5184] ,data[5199:5192] ,data[5207:5200] ,data[5215:5208] ,data[5223:5216] ,data[5415:5408] ,data[5423:5416] ,data[5431:5424] ,data[5439:5432] ,data[5447:5440] ,data[5639:5632] ,data[5647:5640] ,data[5655:5648] ,data[5663:5656] ,data[5671:5664] ,data[5863:5856] ,data[5871:5864] ,data[5879:5872] ,data[5887:5880] ,data[5895:5888] ,data[6087:6080] ,data[6095:6088] ,data[6103:6096] ,data[6111:6104] ,data[6119:6112] };
end
707 :begin
 dPIn = {data[5199:5192] ,data[5207:5200] ,data[5215:5208] ,data[5223:5216] ,data[5231:5224] ,data[5423:5416] ,data[5431:5424] ,data[5439:5432] ,data[5447:5440] ,data[5455:5448] ,data[5647:5640] ,data[5655:5648] ,data[5663:5656] ,data[5671:5664] ,data[5679:5672] ,data[5871:5864] ,data[5879:5872] ,data[5887:5880] ,data[5895:5888] ,data[5903:5896] ,data[6095:6088] ,data[6103:6096] ,data[6111:6104] ,data[6119:6112] ,data[6127:6120] };
end
708 :begin
 dPIn = {data[5207:5200] ,data[5215:5208] ,data[5223:5216] ,data[5231:5224] ,data[5239:5232] ,data[5431:5424] ,data[5439:5432] ,data[5447:5440] ,data[5455:5448] ,data[5463:5456] ,data[5655:5648] ,data[5663:5656] ,data[5671:5664] ,data[5679:5672] ,data[5687:5680] ,data[5879:5872] ,data[5887:5880] ,data[5895:5888] ,data[5903:5896] ,data[5911:5904] ,data[6103:6096] ,data[6111:6104] ,data[6119:6112] ,data[6127:6120] ,data[6135:6128] };
end
709 :begin
 dPIn = {data[5215:5208] ,data[5223:5216] ,data[5231:5224] ,data[5239:5232] ,data[5247:5240] ,data[5439:5432] ,data[5447:5440] ,data[5455:5448] ,data[5463:5456] ,data[5471:5464] ,data[5663:5656] ,data[5671:5664] ,data[5679:5672] ,data[5687:5680] ,data[5695:5688] ,data[5887:5880] ,data[5895:5888] ,data[5903:5896] ,data[5911:5904] ,data[5919:5912] ,data[6111:6104] ,data[6119:6112] ,data[6127:6120] ,data[6135:6128] ,data[6143:6136] };
end
710 :begin
 dPIn = {data[5223:5216] ,data[5231:5224] ,data[5239:5232] ,data[5247:5240] ,data[5255:5248] ,data[5447:5440] ,data[5455:5448] ,data[5463:5456] ,data[5471:5464] ,data[5479:5472] ,data[5671:5664] ,data[5679:5672] ,data[5687:5680] ,data[5695:5688] ,data[5703:5696] ,data[5895:5888] ,data[5903:5896] ,data[5911:5904] ,data[5919:5912] ,data[5927:5920] ,data[6119:6112] ,data[6127:6120] ,data[6135:6128] ,data[6143:6136] ,data[6151:6144] };
end
711 :begin
 dPIn = {data[5231:5224] ,data[5239:5232] ,data[5247:5240] ,data[5255:5248] ,data[5263:5256] ,data[5455:5448] ,data[5463:5456] ,data[5471:5464] ,data[5479:5472] ,data[5487:5480] ,data[5679:5672] ,data[5687:5680] ,data[5695:5688] ,data[5703:5696] ,data[5711:5704] ,data[5903:5896] ,data[5911:5904] ,data[5919:5912] ,data[5927:5920] ,data[5935:5928] ,data[6127:6120] ,data[6135:6128] ,data[6143:6136] ,data[6151:6144] ,data[6159:6152] };
end
712 :begin
 dPIn = {data[5239:5232] ,data[5247:5240] ,data[5255:5248] ,data[5263:5256] ,data[5271:5264] ,data[5463:5456] ,data[5471:5464] ,data[5479:5472] ,data[5487:5480] ,data[5495:5488] ,data[5687:5680] ,data[5695:5688] ,data[5703:5696] ,data[5711:5704] ,data[5719:5712] ,data[5911:5904] ,data[5919:5912] ,data[5927:5920] ,data[5935:5928] ,data[5943:5936] ,data[6135:6128] ,data[6143:6136] ,data[6151:6144] ,data[6159:6152] ,data[6167:6160] };
end
713 :begin
 dPIn = {data[5247:5240] ,data[5255:5248] ,data[5263:5256] ,data[5271:5264] ,data[5279:5272] ,data[5471:5464] ,data[5479:5472] ,data[5487:5480] ,data[5495:5488] ,data[5503:5496] ,data[5695:5688] ,data[5703:5696] ,data[5711:5704] ,data[5719:5712] ,data[5727:5720] ,data[5919:5912] ,data[5927:5920] ,data[5935:5928] ,data[5943:5936] ,data[5951:5944] ,data[6143:6136] ,data[6151:6144] ,data[6159:6152] ,data[6167:6160] ,data[6175:6168] };
end
714 :begin
 dPIn = {data[5255:5248] ,data[5263:5256] ,data[5271:5264] ,data[5279:5272] ,data[5287:5280] ,data[5479:5472] ,data[5487:5480] ,data[5495:5488] ,data[5503:5496] ,data[5511:5504] ,data[5703:5696] ,data[5711:5704] ,data[5719:5712] ,data[5727:5720] ,data[5735:5728] ,data[5927:5920] ,data[5935:5928] ,data[5943:5936] ,data[5951:5944] ,data[5959:5952] ,data[6151:6144] ,data[6159:6152] ,data[6167:6160] ,data[6175:6168] ,data[6183:6176] };
end
715 :begin
 dPIn = {data[5263:5256] ,data[5271:5264] ,data[5279:5272] ,data[5287:5280] ,data[5295:5288] ,data[5487:5480] ,data[5495:5488] ,data[5503:5496] ,data[5511:5504] ,data[5519:5512] ,data[5711:5704] ,data[5719:5712] ,data[5727:5720] ,data[5735:5728] ,data[5743:5736] ,data[5935:5928] ,data[5943:5936] ,data[5951:5944] ,data[5959:5952] ,data[5967:5960] ,data[6159:6152] ,data[6167:6160] ,data[6175:6168] ,data[6183:6176] ,data[6191:6184] };
end
716 :begin
 dPIn = {data[5271:5264] ,data[5279:5272] ,data[5287:5280] ,data[5295:5288] ,data[5303:5296] ,data[5495:5488] ,data[5503:5496] ,data[5511:5504] ,data[5519:5512] ,data[5527:5520] ,data[5719:5712] ,data[5727:5720] ,data[5735:5728] ,data[5743:5736] ,data[5751:5744] ,data[5943:5936] ,data[5951:5944] ,data[5959:5952] ,data[5967:5960] ,data[5975:5968] ,data[6167:6160] ,data[6175:6168] ,data[6183:6176] ,data[6191:6184] ,data[6199:6192] };
end
717 :begin
 dPIn = {data[5279:5272] ,data[5287:5280] ,data[5295:5288] ,data[5303:5296] ,data[5311:5304] ,data[5503:5496] ,data[5511:5504] ,data[5519:5512] ,data[5527:5520] ,data[5535:5528] ,data[5727:5720] ,data[5735:5728] ,data[5743:5736] ,data[5751:5744] ,data[5759:5752] ,data[5951:5944] ,data[5959:5952] ,data[5967:5960] ,data[5975:5968] ,data[5983:5976] ,data[6175:6168] ,data[6183:6176] ,data[6191:6184] ,data[6199:6192] ,data[6207:6200] };
end
718 :begin
 dPIn = {data[5287:5280] ,data[5295:5288] ,data[5303:5296] ,data[5311:5304] ,data[5319:5312] ,data[5511:5504] ,data[5519:5512] ,data[5527:5520] ,data[5535:5528] ,data[5543:5536] ,data[5735:5728] ,data[5743:5736] ,data[5751:5744] ,data[5759:5752] ,data[5767:5760] ,data[5959:5952] ,data[5967:5960] ,data[5975:5968] ,data[5983:5976] ,data[5991:5984] ,data[6183:6176] ,data[6191:6184] ,data[6199:6192] ,data[6207:6200] ,data[6215:6208] };
end
719 :begin
 dPIn = {data[5295:5288] ,data[5303:5296] ,data[5311:5304] ,data[5319:5312] ,data[5327:5320] ,data[5519:5512] ,data[5527:5520] ,data[5535:5528] ,data[5543:5536] ,data[5551:5544] ,data[5743:5736] ,data[5751:5744] ,data[5759:5752] ,data[5767:5760] ,data[5775:5768] ,data[5967:5960] ,data[5975:5968] ,data[5983:5976] ,data[5991:5984] ,data[5999:5992] ,data[6191:6184] ,data[6199:6192] ,data[6207:6200] ,data[6215:6208] ,data[6223:6216] };
end
720 :begin
 dPIn = {data[5303:5296] ,data[5311:5304] ,data[5319:5312] ,data[5327:5320] ,data[5335:5328] ,data[5527:5520] ,data[5535:5528] ,data[5543:5536] ,data[5551:5544] ,data[5559:5552] ,data[5751:5744] ,data[5759:5752] ,data[5767:5760] ,data[5775:5768] ,data[5783:5776] ,data[5975:5968] ,data[5983:5976] ,data[5991:5984] ,data[5999:5992] ,data[6007:6000] ,data[6199:6192] ,data[6207:6200] ,data[6215:6208] ,data[6223:6216] ,data[6231:6224] };
end
721 :begin
 dPIn = {data[5311:5304] ,data[5319:5312] ,data[5327:5320] ,data[5335:5328] ,data[5343:5336] ,data[5535:5528] ,data[5543:5536] ,data[5551:5544] ,data[5559:5552] ,data[5567:5560] ,data[5759:5752] ,data[5767:5760] ,data[5775:5768] ,data[5783:5776] ,data[5791:5784] ,data[5983:5976] ,data[5991:5984] ,data[5999:5992] ,data[6007:6000] ,data[6015:6008] ,data[6207:6200] ,data[6215:6208] ,data[6223:6216] ,data[6231:6224] ,data[6239:6232] };
end
722 :begin
 dPIn = {data[5319:5312] ,data[5327:5320] ,data[5335:5328] ,data[5343:5336] ,data[5351:5344] ,data[5543:5536] ,data[5551:5544] ,data[5559:5552] ,data[5567:5560] ,data[5575:5568] ,data[5767:5760] ,data[5775:5768] ,data[5783:5776] ,data[5791:5784] ,data[5799:5792] ,data[5991:5984] ,data[5999:5992] ,data[6007:6000] ,data[6015:6008] ,data[6023:6016] ,data[6215:6208] ,data[6223:6216] ,data[6231:6224] ,data[6239:6232] ,data[6247:6240] };
end
723 :begin
 dPIn = {data[5327:5320] ,data[5335:5328] ,data[5343:5336] ,data[5351:5344] ,data[5359:5352] ,data[5551:5544] ,data[5559:5552] ,data[5567:5560] ,data[5575:5568] ,data[5583:5576] ,data[5775:5768] ,data[5783:5776] ,data[5791:5784] ,data[5799:5792] ,data[5807:5800] ,data[5999:5992] ,data[6007:6000] ,data[6015:6008] ,data[6023:6016] ,data[6031:6024] ,data[6223:6216] ,data[6231:6224] ,data[6239:6232] ,data[6247:6240] ,data[6255:6248] };
end
724 :begin
 dPIn = {data[5335:5328] ,data[5343:5336] ,data[5351:5344] ,data[5359:5352] ,data[5367:5360] ,data[5559:5552] ,data[5567:5560] ,data[5575:5568] ,data[5583:5576] ,data[5591:5584] ,data[5783:5776] ,data[5791:5784] ,data[5799:5792] ,data[5807:5800] ,data[5815:5808] ,data[6007:6000] ,data[6015:6008] ,data[6023:6016] ,data[6031:6024] ,data[6039:6032] ,data[6231:6224] ,data[6239:6232] ,data[6247:6240] ,data[6255:6248] ,data[6263:6256] };
end
725 :begin
 dPIn = {data[5343:5336] ,data[5351:5344] ,data[5359:5352] ,data[5367:5360] ,data[5375:5368] ,data[5567:5560] ,data[5575:5568] ,data[5583:5576] ,data[5591:5584] ,data[5599:5592] ,data[5791:5784] ,data[5799:5792] ,data[5807:5800] ,data[5815:5808] ,data[5823:5816] ,data[6015:6008] ,data[6023:6016] ,data[6031:6024] ,data[6039:6032] ,data[6047:6040] ,data[6239:6232] ,data[6247:6240] ,data[6255:6248] ,data[6263:6256] ,data[6271:6264] };
end
726 :begin
 dPIn = {data[5351:5344] ,data[5359:5352] ,data[5367:5360] ,data[5375:5368] ,0 ,data[5575:5568] ,data[5583:5576] ,data[5591:5584] ,data[5599:5592] ,0 ,data[5799:5792] ,data[5807:5800] ,data[5815:5808] ,data[5823:5816] ,0 ,data[6023:6016] ,data[6031:6024] ,data[6039:6032] ,data[6047:6040] ,0 ,data[6247:6240] ,data[6255:6248] ,data[6263:6256] ,data[6271:6264] ,0 };
end
727 :begin
 dPIn = {data[5359:5352] ,data[5367:5360] ,data[5375:5368] ,0 ,0 ,data[5583:5576] ,data[5591:5584] ,data[5599:5592] ,0 ,0 ,data[5807:5800] ,data[5815:5808] ,data[5823:5816] ,0 ,0 ,data[6031:6024] ,data[6039:6032] ,data[6047:6040] ,0 ,0 ,data[6255:6248] ,data[6263:6256] ,data[6271:6264] ,0 ,0 };
end
728 :begin
 dPIn = {0 ,0 ,data[5383:5376] ,data[5391:5384] ,data[5399:5392] ,0 ,0 ,data[5607:5600] ,data[5615:5608] ,data[5623:5616] ,0 ,0 ,data[5831:5824] ,data[5839:5832] ,data[5847:5840] ,0 ,0 ,data[6055:6048] ,data[6063:6056] ,data[6071:6064] ,0 ,0 ,0 ,0 ,0 };
end
729 :begin
 dPIn = {0 ,data[5383:5376] ,data[5391:5384] ,data[5399:5392] ,data[5407:5400] ,0 ,data[5607:5600] ,data[5615:5608] ,data[5623:5616] ,data[5631:5624] ,0 ,data[5831:5824] ,data[5839:5832] ,data[5847:5840] ,data[5855:5848] ,0 ,data[6055:6048] ,data[6063:6056] ,data[6071:6064] ,data[6079:6072] ,0 ,0 ,0 ,0 ,0 };
end
730 :begin
 dPIn = {data[5383:5376] ,data[5391:5384] ,data[5399:5392] ,data[5407:5400] ,data[5415:5408] ,data[5607:5600] ,data[5615:5608] ,data[5623:5616] ,data[5631:5624] ,data[5639:5632] ,data[5831:5824] ,data[5839:5832] ,data[5847:5840] ,data[5855:5848] ,data[5863:5856] ,data[6055:6048] ,data[6063:6056] ,data[6071:6064] ,data[6079:6072] ,data[6087:6080] ,0 ,0 ,0 ,0 ,0 };
end
731 :begin
 dPIn = {data[5391:5384] ,data[5399:5392] ,data[5407:5400] ,data[5415:5408] ,data[5423:5416] ,data[5615:5608] ,data[5623:5616] ,data[5631:5624] ,data[5639:5632] ,data[5647:5640] ,data[5839:5832] ,data[5847:5840] ,data[5855:5848] ,data[5863:5856] ,data[5871:5864] ,data[6063:6056] ,data[6071:6064] ,data[6079:6072] ,data[6087:6080] ,data[6095:6088] ,0 ,0 ,0 ,0 ,0 };
end
732 :begin
 dPIn = {data[5399:5392] ,data[5407:5400] ,data[5415:5408] ,data[5423:5416] ,data[5431:5424] ,data[5623:5616] ,data[5631:5624] ,data[5639:5632] ,data[5647:5640] ,data[5655:5648] ,data[5847:5840] ,data[5855:5848] ,data[5863:5856] ,data[5871:5864] ,data[5879:5872] ,data[6071:6064] ,data[6079:6072] ,data[6087:6080] ,data[6095:6088] ,data[6103:6096] ,0 ,0 ,0 ,0 ,0 };
end
733 :begin
 dPIn = {data[5407:5400] ,data[5415:5408] ,data[5423:5416] ,data[5431:5424] ,data[5439:5432] ,data[5631:5624] ,data[5639:5632] ,data[5647:5640] ,data[5655:5648] ,data[5663:5656] ,data[5855:5848] ,data[5863:5856] ,data[5871:5864] ,data[5879:5872] ,data[5887:5880] ,data[6079:6072] ,data[6087:6080] ,data[6095:6088] ,data[6103:6096] ,data[6111:6104] ,0 ,0 ,0 ,0 ,0 };
end
734 :begin
 dPIn = {data[5415:5408] ,data[5423:5416] ,data[5431:5424] ,data[5439:5432] ,data[5447:5440] ,data[5639:5632] ,data[5647:5640] ,data[5655:5648] ,data[5663:5656] ,data[5671:5664] ,data[5863:5856] ,data[5871:5864] ,data[5879:5872] ,data[5887:5880] ,data[5895:5888] ,data[6087:6080] ,data[6095:6088] ,data[6103:6096] ,data[6111:6104] ,data[6119:6112] ,0 ,0 ,0 ,0 ,0 };
end
735 :begin
 dPIn = {data[5423:5416] ,data[5431:5424] ,data[5439:5432] ,data[5447:5440] ,data[5455:5448] ,data[5647:5640] ,data[5655:5648] ,data[5663:5656] ,data[5671:5664] ,data[5679:5672] ,data[5871:5864] ,data[5879:5872] ,data[5887:5880] ,data[5895:5888] ,data[5903:5896] ,data[6095:6088] ,data[6103:6096] ,data[6111:6104] ,data[6119:6112] ,data[6127:6120] ,0 ,0 ,0 ,0 ,0 };
end
736 :begin
 dPIn = {data[5431:5424] ,data[5439:5432] ,data[5447:5440] ,data[5455:5448] ,data[5463:5456] ,data[5655:5648] ,data[5663:5656] ,data[5671:5664] ,data[5679:5672] ,data[5687:5680] ,data[5879:5872] ,data[5887:5880] ,data[5895:5888] ,data[5903:5896] ,data[5911:5904] ,data[6103:6096] ,data[6111:6104] ,data[6119:6112] ,data[6127:6120] ,data[6135:6128] ,0 ,0 ,0 ,0 ,0 };
end
737 :begin
 dPIn = {data[5439:5432] ,data[5447:5440] ,data[5455:5448] ,data[5463:5456] ,data[5471:5464] ,data[5663:5656] ,data[5671:5664] ,data[5679:5672] ,data[5687:5680] ,data[5695:5688] ,data[5887:5880] ,data[5895:5888] ,data[5903:5896] ,data[5911:5904] ,data[5919:5912] ,data[6111:6104] ,data[6119:6112] ,data[6127:6120] ,data[6135:6128] ,data[6143:6136] ,0 ,0 ,0 ,0 ,0 };
end
738 :begin
 dPIn = {data[5447:5440] ,data[5455:5448] ,data[5463:5456] ,data[5471:5464] ,data[5479:5472] ,data[5671:5664] ,data[5679:5672] ,data[5687:5680] ,data[5695:5688] ,data[5703:5696] ,data[5895:5888] ,data[5903:5896] ,data[5911:5904] ,data[5919:5912] ,data[5927:5920] ,data[6119:6112] ,data[6127:6120] ,data[6135:6128] ,data[6143:6136] ,data[6151:6144] ,0 ,0 ,0 ,0 ,0 };
end
739 :begin
 dPIn = {data[5455:5448] ,data[5463:5456] ,data[5471:5464] ,data[5479:5472] ,data[5487:5480] ,data[5679:5672] ,data[5687:5680] ,data[5695:5688] ,data[5703:5696] ,data[5711:5704] ,data[5903:5896] ,data[5911:5904] ,data[5919:5912] ,data[5927:5920] ,data[5935:5928] ,data[6127:6120] ,data[6135:6128] ,data[6143:6136] ,data[6151:6144] ,data[6159:6152] ,0 ,0 ,0 ,0 ,0 };
end
740 :begin
 dPIn = {data[5463:5456] ,data[5471:5464] ,data[5479:5472] ,data[5487:5480] ,data[5495:5488] ,data[5687:5680] ,data[5695:5688] ,data[5703:5696] ,data[5711:5704] ,data[5719:5712] ,data[5911:5904] ,data[5919:5912] ,data[5927:5920] ,data[5935:5928] ,data[5943:5936] ,data[6135:6128] ,data[6143:6136] ,data[6151:6144] ,data[6159:6152] ,data[6167:6160] ,0 ,0 ,0 ,0 ,0 };
end
741 :begin
 dPIn = {data[5471:5464] ,data[5479:5472] ,data[5487:5480] ,data[5495:5488] ,data[5503:5496] ,data[5695:5688] ,data[5703:5696] ,data[5711:5704] ,data[5719:5712] ,data[5727:5720] ,data[5919:5912] ,data[5927:5920] ,data[5935:5928] ,data[5943:5936] ,data[5951:5944] ,data[6143:6136] ,data[6151:6144] ,data[6159:6152] ,data[6167:6160] ,data[6175:6168] ,0 ,0 ,0 ,0 ,0 };
end
742 :begin
 dPIn = {data[5479:5472] ,data[5487:5480] ,data[5495:5488] ,data[5503:5496] ,data[5511:5504] ,data[5703:5696] ,data[5711:5704] ,data[5719:5712] ,data[5727:5720] ,data[5735:5728] ,data[5927:5920] ,data[5935:5928] ,data[5943:5936] ,data[5951:5944] ,data[5959:5952] ,data[6151:6144] ,data[6159:6152] ,data[6167:6160] ,data[6175:6168] ,data[6183:6176] ,0 ,0 ,0 ,0 ,0 };
end
743 :begin
 dPIn = {data[5487:5480] ,data[5495:5488] ,data[5503:5496] ,data[5511:5504] ,data[5519:5512] ,data[5711:5704] ,data[5719:5712] ,data[5727:5720] ,data[5735:5728] ,data[5743:5736] ,data[5935:5928] ,data[5943:5936] ,data[5951:5944] ,data[5959:5952] ,data[5967:5960] ,data[6159:6152] ,data[6167:6160] ,data[6175:6168] ,data[6183:6176] ,data[6191:6184] ,0 ,0 ,0 ,0 ,0 };
end
744 :begin
 dPIn = {data[5495:5488] ,data[5503:5496] ,data[5511:5504] ,data[5519:5512] ,data[5527:5520] ,data[5719:5712] ,data[5727:5720] ,data[5735:5728] ,data[5743:5736] ,data[5751:5744] ,data[5943:5936] ,data[5951:5944] ,data[5959:5952] ,data[5967:5960] ,data[5975:5968] ,data[6167:6160] ,data[6175:6168] ,data[6183:6176] ,data[6191:6184] ,data[6199:6192] ,0 ,0 ,0 ,0 ,0 };
end
745 :begin
 dPIn = {data[5503:5496] ,data[5511:5504] ,data[5519:5512] ,data[5527:5520] ,data[5535:5528] ,data[5727:5720] ,data[5735:5728] ,data[5743:5736] ,data[5751:5744] ,data[5759:5752] ,data[5951:5944] ,data[5959:5952] ,data[5967:5960] ,data[5975:5968] ,data[5983:5976] ,data[6175:6168] ,data[6183:6176] ,data[6191:6184] ,data[6199:6192] ,data[6207:6200] ,0 ,0 ,0 ,0 ,0 };
end
746 :begin
 dPIn = {data[5511:5504] ,data[5519:5512] ,data[5527:5520] ,data[5535:5528] ,data[5543:5536] ,data[5735:5728] ,data[5743:5736] ,data[5751:5744] ,data[5759:5752] ,data[5767:5760] ,data[5959:5952] ,data[5967:5960] ,data[5975:5968] ,data[5983:5976] ,data[5991:5984] ,data[6183:6176] ,data[6191:6184] ,data[6199:6192] ,data[6207:6200] ,data[6215:6208] ,0 ,0 ,0 ,0 ,0 };
end
747 :begin
 dPIn = {data[5519:5512] ,data[5527:5520] ,data[5535:5528] ,data[5543:5536] ,data[5551:5544] ,data[5743:5736] ,data[5751:5744] ,data[5759:5752] ,data[5767:5760] ,data[5775:5768] ,data[5967:5960] ,data[5975:5968] ,data[5983:5976] ,data[5991:5984] ,data[5999:5992] ,data[6191:6184] ,data[6199:6192] ,data[6207:6200] ,data[6215:6208] ,data[6223:6216] ,0 ,0 ,0 ,0 ,0 };
end
748 :begin
 dPIn = {data[5527:5520] ,data[5535:5528] ,data[5543:5536] ,data[5551:5544] ,data[5559:5552] ,data[5751:5744] ,data[5759:5752] ,data[5767:5760] ,data[5775:5768] ,data[5783:5776] ,data[5975:5968] ,data[5983:5976] ,data[5991:5984] ,data[5999:5992] ,data[6007:6000] ,data[6199:6192] ,data[6207:6200] ,data[6215:6208] ,data[6223:6216] ,data[6231:6224] ,0 ,0 ,0 ,0 ,0 };
end
749 :begin
 dPIn = {data[5535:5528] ,data[5543:5536] ,data[5551:5544] ,data[5559:5552] ,data[5567:5560] ,data[5759:5752] ,data[5767:5760] ,data[5775:5768] ,data[5783:5776] ,data[5791:5784] ,data[5983:5976] ,data[5991:5984] ,data[5999:5992] ,data[6007:6000] ,data[6015:6008] ,data[6207:6200] ,data[6215:6208] ,data[6223:6216] ,data[6231:6224] ,data[6239:6232] ,0 ,0 ,0 ,0 ,0 };
end
750 :begin
 dPIn = {data[5543:5536] ,data[5551:5544] ,data[5559:5552] ,data[5567:5560] ,data[5575:5568] ,data[5767:5760] ,data[5775:5768] ,data[5783:5776] ,data[5791:5784] ,data[5799:5792] ,data[5991:5984] ,data[5999:5992] ,data[6007:6000] ,data[6015:6008] ,data[6023:6016] ,data[6215:6208] ,data[6223:6216] ,data[6231:6224] ,data[6239:6232] ,data[6247:6240] ,0 ,0 ,0 ,0 ,0 };
end
751 :begin
 dPIn = {data[5551:5544] ,data[5559:5552] ,data[5567:5560] ,data[5575:5568] ,data[5583:5576] ,data[5775:5768] ,data[5783:5776] ,data[5791:5784] ,data[5799:5792] ,data[5807:5800] ,data[5999:5992] ,data[6007:6000] ,data[6015:6008] ,data[6023:6016] ,data[6031:6024] ,data[6223:6216] ,data[6231:6224] ,data[6239:6232] ,data[6247:6240] ,data[6255:6248] ,0 ,0 ,0 ,0 ,0 };
end
752 :begin
 dPIn = {data[5559:5552] ,data[5567:5560] ,data[5575:5568] ,data[5583:5576] ,data[5591:5584] ,data[5783:5776] ,data[5791:5784] ,data[5799:5792] ,data[5807:5800] ,data[5815:5808] ,data[6007:6000] ,data[6015:6008] ,data[6023:6016] ,data[6031:6024] ,data[6039:6032] ,data[6231:6224] ,data[6239:6232] ,data[6247:6240] ,data[6255:6248] ,data[6263:6256] ,0 ,0 ,0 ,0 ,0 };
end
753 :begin
 dPIn = {data[5567:5560] ,data[5575:5568] ,data[5583:5576] ,data[5591:5584] ,data[5599:5592] ,data[5791:5784] ,data[5799:5792] ,data[5807:5800] ,data[5815:5808] ,data[5823:5816] ,data[6015:6008] ,data[6023:6016] ,data[6031:6024] ,data[6039:6032] ,data[6047:6040] ,data[6239:6232] ,data[6247:6240] ,data[6255:6248] ,data[6263:6256] ,data[6271:6264] ,0 ,0 ,0 ,0 ,0 };
end
754 :begin
 dPIn = {data[5575:5568] ,data[5583:5576] ,data[5591:5584] ,data[5599:5592] ,0 ,data[5799:5792] ,data[5807:5800] ,data[5815:5808] ,data[5823:5816] ,0 ,data[6023:6016] ,data[6031:6024] ,data[6039:6032] ,data[6047:6040] ,0 ,data[6247:6240] ,data[6255:6248] ,data[6263:6256] ,data[6271:6264] ,0 ,0 ,0 ,0 ,0 ,0 };
end
755 :begin
 dPIn = {data[5583:5576] ,data[5591:5584] ,data[5599:5592] ,0 ,0 ,data[5807:5800] ,data[5815:5808] ,data[5823:5816] ,0 ,0 ,data[6031:6024] ,data[6039:6032] ,data[6047:6040] ,0 ,0 ,data[6255:6248] ,data[6263:6256] ,data[6271:6264] ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
756 :begin
 dPIn = {0 ,0 ,data[5607:5600] ,data[5615:5608] ,data[5623:5616] ,0 ,0 ,data[5831:5824] ,data[5839:5832] ,data[5847:5840] ,0 ,0 ,data[6055:6048] ,data[6063:6056] ,data[6071:6064] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
757 :begin
 dPIn = {0 ,data[5607:5600] ,data[5615:5608] ,data[5623:5616] ,data[5631:5624] ,0 ,data[5831:5824] ,data[5839:5832] ,data[5847:5840] ,data[5855:5848] ,0 ,data[6055:6048] ,data[6063:6056] ,data[6071:6064] ,data[6079:6072] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
758 :begin
 dPIn = {data[5607:5600] ,data[5615:5608] ,data[5623:5616] ,data[5631:5624] ,data[5639:5632] ,data[5831:5824] ,data[5839:5832] ,data[5847:5840] ,data[5855:5848] ,data[5863:5856] ,data[6055:6048] ,data[6063:6056] ,data[6071:6064] ,data[6079:6072] ,data[6087:6080] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
759 :begin
 dPIn = {data[5615:5608] ,data[5623:5616] ,data[5631:5624] ,data[5639:5632] ,data[5647:5640] ,data[5839:5832] ,data[5847:5840] ,data[5855:5848] ,data[5863:5856] ,data[5871:5864] ,data[6063:6056] ,data[6071:6064] ,data[6079:6072] ,data[6087:6080] ,data[6095:6088] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
760 :begin
 dPIn = {data[5623:5616] ,data[5631:5624] ,data[5639:5632] ,data[5647:5640] ,data[5655:5648] ,data[5847:5840] ,data[5855:5848] ,data[5863:5856] ,data[5871:5864] ,data[5879:5872] ,data[6071:6064] ,data[6079:6072] ,data[6087:6080] ,data[6095:6088] ,data[6103:6096] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
761 :begin
 dPIn = {data[5631:5624] ,data[5639:5632] ,data[5647:5640] ,data[5655:5648] ,data[5663:5656] ,data[5855:5848] ,data[5863:5856] ,data[5871:5864] ,data[5879:5872] ,data[5887:5880] ,data[6079:6072] ,data[6087:6080] ,data[6095:6088] ,data[6103:6096] ,data[6111:6104] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
762 :begin
 dPIn = {data[5639:5632] ,data[5647:5640] ,data[5655:5648] ,data[5663:5656] ,data[5671:5664] ,data[5863:5856] ,data[5871:5864] ,data[5879:5872] ,data[5887:5880] ,data[5895:5888] ,data[6087:6080] ,data[6095:6088] ,data[6103:6096] ,data[6111:6104] ,data[6119:6112] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
763 :begin
 dPIn = {data[5647:5640] ,data[5655:5648] ,data[5663:5656] ,data[5671:5664] ,data[5679:5672] ,data[5871:5864] ,data[5879:5872] ,data[5887:5880] ,data[5895:5888] ,data[5903:5896] ,data[6095:6088] ,data[6103:6096] ,data[6111:6104] ,data[6119:6112] ,data[6127:6120] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
764 :begin
 dPIn = {data[5655:5648] ,data[5663:5656] ,data[5671:5664] ,data[5679:5672] ,data[5687:5680] ,data[5879:5872] ,data[5887:5880] ,data[5895:5888] ,data[5903:5896] ,data[5911:5904] ,data[6103:6096] ,data[6111:6104] ,data[6119:6112] ,data[6127:6120] ,data[6135:6128] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
765 :begin
 dPIn = {data[5663:5656] ,data[5671:5664] ,data[5679:5672] ,data[5687:5680] ,data[5695:5688] ,data[5887:5880] ,data[5895:5888] ,data[5903:5896] ,data[5911:5904] ,data[5919:5912] ,data[6111:6104] ,data[6119:6112] ,data[6127:6120] ,data[6135:6128] ,data[6143:6136] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
766 :begin
 dPIn = {data[5671:5664] ,data[5679:5672] ,data[5687:5680] ,data[5695:5688] ,data[5703:5696] ,data[5895:5888] ,data[5903:5896] ,data[5911:5904] ,data[5919:5912] ,data[5927:5920] ,data[6119:6112] ,data[6127:6120] ,data[6135:6128] ,data[6143:6136] ,data[6151:6144] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
767 :begin
 dPIn = {data[5679:5672] ,data[5687:5680] ,data[5695:5688] ,data[5703:5696] ,data[5711:5704] ,data[5903:5896] ,data[5911:5904] ,data[5919:5912] ,data[5927:5920] ,data[5935:5928] ,data[6127:6120] ,data[6135:6128] ,data[6143:6136] ,data[6151:6144] ,data[6159:6152] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
768 :begin
 dPIn = {data[5687:5680] ,data[5695:5688] ,data[5703:5696] ,data[5711:5704] ,data[5719:5712] ,data[5911:5904] ,data[5919:5912] ,data[5927:5920] ,data[5935:5928] ,data[5943:5936] ,data[6135:6128] ,data[6143:6136] ,data[6151:6144] ,data[6159:6152] ,data[6167:6160] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
769 :begin
 dPIn = {data[5695:5688] ,data[5703:5696] ,data[5711:5704] ,data[5719:5712] ,data[5727:5720] ,data[5919:5912] ,data[5927:5920] ,data[5935:5928] ,data[5943:5936] ,data[5951:5944] ,data[6143:6136] ,data[6151:6144] ,data[6159:6152] ,data[6167:6160] ,data[6175:6168] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
770 :begin
 dPIn = {data[5703:5696] ,data[5711:5704] ,data[5719:5712] ,data[5727:5720] ,data[5735:5728] ,data[5927:5920] ,data[5935:5928] ,data[5943:5936] ,data[5951:5944] ,data[5959:5952] ,data[6151:6144] ,data[6159:6152] ,data[6167:6160] ,data[6175:6168] ,data[6183:6176] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
771 :begin
 dPIn = {data[5711:5704] ,data[5719:5712] ,data[5727:5720] ,data[5735:5728] ,data[5743:5736] ,data[5935:5928] ,data[5943:5936] ,data[5951:5944] ,data[5959:5952] ,data[5967:5960] ,data[6159:6152] ,data[6167:6160] ,data[6175:6168] ,data[6183:6176] ,data[6191:6184] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
772 :begin
 dPIn = {data[5719:5712] ,data[5727:5720] ,data[5735:5728] ,data[5743:5736] ,data[5751:5744] ,data[5943:5936] ,data[5951:5944] ,data[5959:5952] ,data[5967:5960] ,data[5975:5968] ,data[6167:6160] ,data[6175:6168] ,data[6183:6176] ,data[6191:6184] ,data[6199:6192] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
773 :begin
 dPIn = {data[5727:5720] ,data[5735:5728] ,data[5743:5736] ,data[5751:5744] ,data[5759:5752] ,data[5951:5944] ,data[5959:5952] ,data[5967:5960] ,data[5975:5968] ,data[5983:5976] ,data[6175:6168] ,data[6183:6176] ,data[6191:6184] ,data[6199:6192] ,data[6207:6200] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
774 :begin
 dPIn = {data[5735:5728] ,data[5743:5736] ,data[5751:5744] ,data[5759:5752] ,data[5767:5760] ,data[5959:5952] ,data[5967:5960] ,data[5975:5968] ,data[5983:5976] ,data[5991:5984] ,data[6183:6176] ,data[6191:6184] ,data[6199:6192] ,data[6207:6200] ,data[6215:6208] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
775 :begin
 dPIn = {data[5743:5736] ,data[5751:5744] ,data[5759:5752] ,data[5767:5760] ,data[5775:5768] ,data[5967:5960] ,data[5975:5968] ,data[5983:5976] ,data[5991:5984] ,data[5999:5992] ,data[6191:6184] ,data[6199:6192] ,data[6207:6200] ,data[6215:6208] ,data[6223:6216] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
776 :begin
 dPIn = {data[5751:5744] ,data[5759:5752] ,data[5767:5760] ,data[5775:5768] ,data[5783:5776] ,data[5975:5968] ,data[5983:5976] ,data[5991:5984] ,data[5999:5992] ,data[6007:6000] ,data[6199:6192] ,data[6207:6200] ,data[6215:6208] ,data[6223:6216] ,data[6231:6224] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
777 :begin
 dPIn = {data[5759:5752] ,data[5767:5760] ,data[5775:5768] ,data[5783:5776] ,data[5791:5784] ,data[5983:5976] ,data[5991:5984] ,data[5999:5992] ,data[6007:6000] ,data[6015:6008] ,data[6207:6200] ,data[6215:6208] ,data[6223:6216] ,data[6231:6224] ,data[6239:6232] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
778 :begin
 dPIn = {data[5767:5760] ,data[5775:5768] ,data[5783:5776] ,data[5791:5784] ,data[5799:5792] ,data[5991:5984] ,data[5999:5992] ,data[6007:6000] ,data[6015:6008] ,data[6023:6016] ,data[6215:6208] ,data[6223:6216] ,data[6231:6224] ,data[6239:6232] ,data[6247:6240] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
779 :begin
 dPIn = {data[5775:5768] ,data[5783:5776] ,data[5791:5784] ,data[5799:5792] ,data[5807:5800] ,data[5999:5992] ,data[6007:6000] ,data[6015:6008] ,data[6023:6016] ,data[6031:6024] ,data[6223:6216] ,data[6231:6224] ,data[6239:6232] ,data[6247:6240] ,data[6255:6248] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
780 :begin
 dPIn = {data[5783:5776] ,data[5791:5784] ,data[5799:5792] ,data[5807:5800] ,data[5815:5808] ,data[6007:6000] ,data[6015:6008] ,data[6023:6016] ,data[6031:6024] ,data[6039:6032] ,data[6231:6224] ,data[6239:6232] ,data[6247:6240] ,data[6255:6248] ,data[6263:6256] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
781 :begin
 dPIn = {data[5791:5784] ,data[5799:5792] ,data[5807:5800] ,data[5815:5808] ,data[5823:5816] ,data[6015:6008] ,data[6023:6016] ,data[6031:6024] ,data[6039:6032] ,data[6047:6040] ,data[6239:6232] ,data[6247:6240] ,data[6255:6248] ,data[6263:6256] ,data[6271:6264] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
782 :begin
 dPIn = {data[5799:5792] ,data[5807:5800] ,data[5815:5808] ,data[5823:5816] ,0 ,data[6023:6016] ,data[6031:6024] ,data[6039:6032] ,data[6047:6040] ,0 ,data[6247:6240] ,data[6255:6248] ,data[6263:6256] ,data[6271:6264] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
783 :begin
 dPIn = {data[5807:5800] ,data[5815:5808] ,data[5823:5816] ,0 ,0 ,data[6031:6024] ,data[6039:6032] ,data[6047:6040] ,0 ,0 ,data[6255:6248] ,data[6263:6256] ,data[6271:6264] ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 ,0 };
end
endcase

end
endmodule

